`include "accel_src/mem_Accel_B.v"

module Htif(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    output io_cpu_0_reset,
    output io_cpu_0_id,
    input  io_cpu_0_csr_req_ready,
    output io_cpu_0_csr_req_valid,
    output io_cpu_0_csr_req_bits_rw,
    output[11:0] io_cpu_0_csr_req_bits_addr,
    output[63:0] io_cpu_0_csr_req_bits_data,
    output io_cpu_0_csr_resp_ready,
    input  io_cpu_0_csr_resp_valid,
    input [63:0] io_cpu_0_csr_resp_bits,
    input  io_cpu_0_debug_stats_csr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[5:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits
);

  wire[63:0] csr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  reg [2:0] state;
  wire[2:0] T210;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T211;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T212;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire[39:0] T50;
  wire[39:0] T51;
  wire T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T213;
  wire[14:0] T57;
  wire[14:0] T58;
  wire[14:0] T59;
  wire T60;
  wire T61;
  wire[3:0] next_cmd;
  wire T62;
  wire[12:0] rx_word_count;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire rx_done;
  wire T67;
  wire T68;
  wire T69;
  wire[2:0] T70;
  wire T71;
  wire[12:0] T214;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire rx_word_done;
  wire T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire cnt_done;
  wire T80;
  reg [1:0] cnt;
  wire[1:0] T215;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  reg [8:0] pos;
  wire[8:0] T94;
  wire[8:0] T95;
  wire[8:0] T96;
  wire[8:0] T97;
  wire[8:0] T98;
  wire[8:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[2:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire tx_done;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire[12:0] T216;
  wire T120;
  wire T121;
  wire[1:0] tx_subword_count;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[11:0] csr_addr;
  wire T126;
  wire T127;
  wire[1:0] csr_coreid;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[63:0] T135;
  wire[63:0] T136;
  wire T137;
  wire T138;
  wire[2:0] T139;
  wire[63:0] T140;
  wire T141;
  wire[2:0] T142;
  wire[2:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[127:0] T150;
  wire[127:0] T151;
  wire[127:0] T152;
  wire[127:0] mem_req_data;
  wire[63:0] T153;
  wire[2:0] T154;
  wire[63:0] T155;
  wire[2:0] T156;
  wire T157;
  wire[16:0] T158;
  wire[16:0] T159;
  wire[16:0] T160;
  wire[16:0] T161;
  wire[15:0] T162;
  wire[2:0] T163;
  wire[2:0] T164;
  wire[2:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[5:0] T172;
  wire[5:0] T173;
  wire[5:0] T174;
  wire[25:0] T175;
  wire[25:0] T176;
  wire[25:0] T217;
  wire[36:0] init_addr;
  wire[39:0] T177;
  wire[25:0] T178;
  wire[25:0] T218;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg  R187;
  wire T219;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire[15:0] T220;
  wire[63:0] T192;
  wire[5:0] T193;
  wire[1:0] T194;
  wire[63:0] tx_data;
  wire[63:0] T195;
  wire[63:0] T196;
  reg [63:0] csrReadData;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T199;
  wire[63:0] T221;
  wire T200;
  wire T201;
  wire T202;
  wire[63:0] tx_header;
  wire[15:0] T203;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T204;
  reg [7:0] seqno;
  wire[7:0] T205;
  wire[7:0] T206;
  wire T207;
  wire T208;
  wire T209;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    state = {1{$random}};
    cmd = {1{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    rx_shifter = {2{$random}};
    addr = {2{$random}};
    tx_count = {1{$random}};
    cnt = {1{$random}};
    pos = {1{$random}};
    R187 = {1{$random}};
    csrReadData = {2{$random}};
    seqno = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign io_cpu_0_id = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_scr_resp_ready = 1'h1;
  assign io_scr_req_bits_data = csr_wdata;
  assign csr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_data[7'h7f:7'h40];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 3'h5;
  assign T210 = reset ? 3'h0 : T4;
  assign T4 = T132 ? 3'h7 : T5;
  assign T5 = T131 ? 3'h2 : T6;
  assign T6 = T129 ? 3'h7 : T7;
  assign T7 = T124 ? 3'h7 : T8;
  assign T8 = T123 ? 3'h2 : T9;
  assign T9 = T113 ? T109 : T10;
  assign T10 = T107 ? T103 : T11;
  assign T11 = T101 ? T91 : T12;
  assign T12 = T89 ? 3'h5 : T13;
  assign T13 = T79 ? 3'h6 : T14;
  assign T14 = T66 ? T15 : state;
  assign T15 = T65 ? 3'h3 : T16;
  assign T16 = T64 ? 3'h4 : T17;
  assign T17 = T18 ? 3'h1 : 3'h7;
  assign T18 = T63 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T62 ? next_cmd : cmd;
  assign T20 = T21 ? next_cmd : cmd;
  assign T21 = T61 & T22;
  assign T22 = rx_count == 15'h3;
  assign T211 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T61 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T113 & T27;
  assign T27 = tx_word_count == T212;
  assign T212 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T61 ? rx_shifter_in : rx_shifter;
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T54 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T52 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T107 ? T51 : T47;
  assign T47 = T101 ? T50 : T48;
  assign T48 = T21 ? T49 : addr;
  assign T49 = rx_shifter_in[6'h3f:5'h18];
  assign T50 = addr + 40'h8;
  assign T51 = addr + 40'h8;
  assign T52 = T53 != 3'h0;
  assign T53 = size[2'h2:1'h0];
  assign T54 = T56 | T55;
  assign T55 = cmd == 4'h1;
  assign T56 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T213 = reset ? 15'h0 : T57;
  assign T57 = T26 ? 15'h0 : T58;
  assign T58 = T60 ? T59 : tx_count;
  assign T59 = tx_count + 15'h1;
  assign T60 = io_host_out_valid & io_host_out_ready;
  assign T61 = io_host_in_valid & io_host_in_ready;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign T62 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T63 = rx_cmd == 4'h2;
  assign T64 = rx_cmd == 4'h1;
  assign T65 = rx_cmd == 4'h0;
  assign T66 = T78 & rx_done;
  assign rx_done = rx_word_done & T67;
  assign T67 = T75 ? T72 : T68;
  assign T68 = T71 | T69;
  assign T69 = T70 == 3'h0;
  assign T70 = rx_word_count[2'h2:1'h0];
  assign T71 = rx_word_count == T214;
  assign T214 = {1'h0, size};
  assign T72 = T74 & T73;
  assign T73 = next_cmd != 4'h3;
  assign T74 = next_cmd != 4'h1;
  assign T75 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T76;
  assign T76 = T77 == 2'h3;
  assign T77 = rx_count[1'h1:1'h0];
  assign T78 = state == 3'h0;
  assign T79 = T88 & cnt_done;
  assign cnt_done = T83 & T80;
  assign T80 = cnt == 2'h3;
  assign T215 = reset ? 2'h0 : T81;
  assign T81 = T83 ? T82 : cnt;
  assign T82 = cnt + 2'h1;
  assign T83 = T86 | T84;
  assign T84 = T85 & io_mem_grant_valid;
  assign T85 = state == 3'h5;
  assign T86 = T87 & io_mem_acquire_ready;
  assign T87 = state == 3'h4;
  assign T88 = state == 3'h4;
  assign T89 = T90 & io_mem_acquire_ready;
  assign T90 = state == 3'h3;
  assign T91 = T92 ? 3'h7 : 3'h0;
  assign T92 = T100 | T93;
  assign T93 = pos == 9'h1;
  assign T94 = T107 ? T99 : T95;
  assign T95 = T101 ? T98 : T96;
  assign T96 = T21 ? T97 : pos;
  assign T97 = rx_shifter_in[4'hf:3'h7];
  assign T98 = pos - 9'h1;
  assign T99 = pos - 9'h1;
  assign T100 = cmd == 4'h0;
  assign T101 = T102 & io_mem_grant_valid;
  assign T102 = state == 3'h6;
  assign T103 = T104 ? 3'h7 : 3'h0;
  assign T104 = T106 | T105;
  assign T105 = pos == 9'h1;
  assign T106 = cmd == 4'h0;
  assign T107 = T108 & cnt_done;
  assign T108 = state == 3'h5;
  assign T109 = T110 ? 3'h3 : 3'h0;
  assign T110 = T112 & T111;
  assign T111 = pos != 9'h0;
  assign T112 = cmd == 4'h0;
  assign T113 = T122 & tx_done;
  assign tx_done = T120 & T114;
  assign T114 = T119 | T115;
  assign T115 = T118 & T116;
  assign T116 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T117 - 3'h1;
  assign T117 = tx_word_count[2'h2:1'h0];
  assign T118 = 13'h0 < tx_word_count;
  assign T119 = tx_word_count == T216;
  assign T216 = {1'h0, tx_size};
  assign T120 = io_host_out_ready & T121;
  assign T121 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T122 = state == 3'h7;
  assign T123 = io_cpu_0_csr_req_ready & io_cpu_0_csr_req_valid;
  assign T124 = T126 & T125;
  assign T125 = csr_addr == 12'h782;
  assign csr_addr = addr[4'hb:1'h0];
  assign T126 = T128 & T127;
  assign T127 = csr_coreid == 2'h0;
  assign csr_coreid = addr[5'h15:5'h14];
  assign T128 = state == 3'h1;
  assign T129 = T130 & io_cpu_0_csr_resp_valid;
  assign T130 = state == 3'h2;
  assign T131 = io_scr_req_ready & io_scr_req_valid;
  assign T132 = T133 & io_scr_resp_valid;
  assign T133 = state == 3'h2;
  assign T134 = {io_mem_grant_bits_addr_beat, 1'h1};
  assign T136 = io_mem_grant_bits_data[6'h3f:1'h0];
  assign T137 = T138 & io_mem_grant_valid;
  assign T138 = state == 3'h5;
  assign T139 = {io_mem_grant_bits_addr_beat, 1'h0};
  assign T141 = rx_word_done & io_host_in_ready;
  assign T142 = T143 - 3'h1;
  assign T143 = rx_word_count[2'h2:1'h0];
  assign io_scr_req_bits_addr = T144;
  assign T144 = T145;
  assign T145 = addr[3'h5:1'h0];
  assign io_scr_req_bits_rw = T146;
  assign T146 = cmd == 4'h3;
  assign io_scr_req_valid = T147;
  assign T147 = T149 & T148;
  assign T148 = csr_coreid == 2'h3;
  assign T149 = state == 3'h1;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_data = T150;
  assign T150 = T157 ? T152 : T151;
  assign T151 = 128'h0;
  assign T152 = mem_req_data;
  assign mem_req_data = {T155, T153};
  assign T153 = packet_ram[T154];
  assign T154 = {cnt, 1'h0};
  assign T155 = packet_ram[T156];
  assign T156 = {cnt, 1'h1};
  assign T157 = cmd == 4'h1;
  assign io_mem_acquire_bits_union = T158;
  assign T158 = T157 ? T160 : T159;
  assign T159 = 17'h1c1;
  assign T160 = T161;
  assign T161 = {T162, 1'h1};
  assign T162 = 16'hffff;
  assign io_mem_acquire_bits_a_type = T163;
  assign T163 = T157 ? T165 : T164;
  assign T164 = 3'h1;
  assign T165 = 3'h3;
  assign io_mem_acquire_bits_is_builtin_type = T166;
  assign T166 = T157 ? T168 : T167;
  assign T167 = 1'h1;
  assign T168 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T169;
  assign T169 = T157 ? T171 : T170;
  assign T170 = 2'h0;
  assign T171 = cnt;
  assign io_mem_acquire_bits_client_xact_id = T172;
  assign T172 = T157 ? T174 : T173;
  assign T173 = 6'h0;
  assign T174 = 6'h0;
  assign io_mem_acquire_bits_addr_block = T175;
  assign T175 = T157 ? T178 : T176;
  assign T176 = T217;
  assign T217 = init_addr[5'h19:1'h0];
  assign init_addr = T177 >> 2'h3;
  assign T177 = addr;
  assign T178 = T218;
  assign T218 = init_addr[5'h19:1'h0];
  assign io_mem_acquire_valid = T179;
  assign T179 = T181 | T180;
  assign T180 = state == 3'h4;
  assign T181 = state == 3'h3;
  assign io_cpu_0_csr_resp_ready = 1'h1;
  assign io_cpu_0_csr_req_bits_data = csr_wdata;
  assign io_cpu_0_csr_req_bits_addr = csr_addr;
  assign io_cpu_0_csr_req_bits_rw = T182;
  assign T182 = cmd == 4'h3;
  assign io_cpu_0_csr_req_valid = T183;
  assign T183 = T185 & T184;
  assign T184 = csr_addr != 12'h782;
  assign T185 = T186 & T127;
  assign T186 = state == 3'h1;
  assign io_cpu_0_reset = R187;
  assign T219 = reset ? 1'h1 : T188;
  assign T188 = T190 ? T189 : R187;
  assign T189 = csr_wdata[1'h0];
  assign T190 = T124 & T191;
  assign T191 = cmd == 4'h3;
  assign io_host_debug_stats_csr = io_cpu_0_debug_stats_csr;
  assign io_host_out_bits = T220;
  assign T220 = T192[4'hf:1'h0];
  assign T192 = tx_data >> T193;
  assign T193 = {T194, 4'h0};
  assign T194 = tx_count[1'h1:1'h0];
  assign tx_data = T207 ? tx_header : T195;
  assign T195 = T200 ? csrReadData : T196;
  assign T196 = packet_ram[packet_ram_raddr];
  assign T197 = T132 ? io_scr_resp_bits : T198;
  assign T198 = T129 ? io_cpu_0_csr_resp_bits : T199;
  assign T199 = T124 ? T221 : csrReadData;
  assign T221 = {63'h0, R187};
  assign T200 = T202 | T201;
  assign T201 = cmd == 4'h3;
  assign T202 = cmd == 4'h2;
  assign tx_header = {T204, T203};
  assign T203 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T204 = {addr, seqno};
  assign T205 = T21 ? T206 : seqno;
  assign T206 = rx_shifter_in[5'h17:5'h10];
  assign T207 = tx_word_count == 13'h0;
  assign io_host_out_valid = T208;
  assign T208 = state == 3'h7;
  assign io_host_in_ready = T209;
  assign T209 = state == 3'h0;

  always @(posedge clk) begin
    if (T2)
      packet_ram[T134] <= T1;
    if(reset) begin
      state <= 3'h0;
    end else if(T132) begin
      state <= 3'h7;
    end else if(T131) begin
      state <= 3'h2;
    end else if(T129) begin
      state <= 3'h7;
    end else if(T124) begin
      state <= 3'h7;
    end else if(T123) begin
      state <= 3'h2;
    end else if(T113) begin
      state <= T109;
    end else if(T107) begin
      state <= T103;
    end else if(T101) begin
      state <= T91;
    end else if(T89) begin
      state <= 3'h5;
    end else if(T79) begin
      state <= 3'h6;
    end else if(T66) begin
      state <= T15;
    end
    if(T21) begin
      cmd <= next_cmd;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T61) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T61) begin
      rx_shifter <= rx_shifter_in;
    end
    if(T107) begin
      addr <= T51;
    end else if(T101) begin
      addr <= T50;
    end else if(T21) begin
      addr <= T49;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T60) begin
      tx_count <= T59;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T83) begin
      cnt <= T82;
    end
    if(T107) begin
      pos <= T99;
    end else if(T101) begin
      pos <= T98;
    end else if(T21) begin
      pos <= T97;
    end
    if (T137)
      packet_ram[T139] <= T136;
    if (T141)
      packet_ram[T142] <= rx_shifter_in;
    if(reset) begin
      R187 <= 1'h1;
    end else if(T190) begin
      R187 <= T189;
    end
    if(T132) begin
      csrReadData <= io_scr_resp_bits;
    end else if(T129) begin
      csrReadData <= io_cpu_0_csr_resp_bits;
    end else if(T124) begin
      csrReadData <= T221;
    end
    if(T21) begin
      seqno <= T206;
    end
  end
endmodule

module ClientTileLinkIOWrapper_0(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [5:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[5:0] io_in_grant_bits_client_xact_id,
    output[3:0] io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[5:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [5:0] io_out_grant_bits_client_xact_id,
    input [3:0] io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[5:0] io_out_release_bits_client_xact_id
    //output io_out_release_bits_voluntary
    //output[2:0] io_out_release_bits_r_type
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module FinishQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [3:0] io_enq_bits_fin_manager_xact_id,
    input [2:0] io_enq_bits_dst,
    input  io_deq_ready,
    output io_deq_valid,
    output[3:0] io_deq_bits_fin_manager_xact_id,
    output[2:0] io_deq_bits_dst,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[6:0] T11;
  reg [6:0] ram [1:0];
  wire[6:0] T12;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[3:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_dst = T10;
  assign T10 = T11[2'h2:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_fin_manager_xact_id, io_enq_bits_dst};
  assign io_deq_bits_fin_manager_xact_id = T15;
  assign T15 = T11[3'h6:2'h3];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module FinishUnit_0(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [2:0] io_grant_bits_header_src,
    input [2:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [5:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[5:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[2:0] io_finish_bits_header_src,
    output[2:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[2:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 3'h0;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [5:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[5:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [5:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[2:0] io_network_acquire_bits_header_src,
    output[2:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[5:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [2:0] io_network_grant_bits_header_src,
    input [2:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [5:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[2:0] io_network_finish_bits_header_src,
    output[2:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [2:0] io_network_probe_bits_header_src,
    input [2:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[2:0] io_network_release_bits_header_src,
    output[2:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[5:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[5:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[2:0] rel_with_header_bits_header_dst;
  wire[2:0] T8;
  wire T0;
  wire T1;
  wire[25:0] T2;
  wire[2:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[5:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[2:0] acq_with_header_bits_header_dst;
  wire[2:0] T9;
  wire T3;
  wire T4;
  wire[25:0] T5;
  wire[2:0] acq_with_header_bits_header_src;
  wire T6;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T7;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[5:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[2:0] finisher_io_finish_bits_header_src;
  wire[2:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = T8;
  assign T8 = {2'h0, T0};
  assign T0 = T1 == 1'h0;
  assign T1 = T2 < 26'h1000000;
  assign T2 = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 3'h0;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = T9;
  assign T9 = {2'h0, T3};
  assign T3 = T4 == 1'h0;
  assign T4 = T5 < 26'h1000000;
  assign T5 = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 3'h0;
  assign io_network_acquire_valid = T6;
  assign T6 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T7;
  assign T7 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_0 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [5:0] io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input  io_enq_bits_payload_is_builtin_type,
    input [2:0] io_enq_bits_payload_a_type,
    input [16:0] io_enq_bits_payload_union,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[5:0] io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output io_deq_bits_payload_is_builtin_type,
    output[2:0] io_deq_bits_payload_a_type,
    output[16:0] io_deq_bits_payload_union,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T33;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T34;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T35;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[188:0] T11;
  reg [188:0] ram [1:0];
  wire[188:0] T12;
  wire[188:0] T13;
  wire[188:0] T14;
  wire[150:0] T15;
  wire[147:0] T16;
  wire[144:0] T17;
  wire[2:0] T18;
  wire[37:0] T19;
  wire[31:0] T20;
  wire[5:0] T21;
  wire[16:0] T22;
  wire[2:0] T23;
  wire T24;
  wire[1:0] T25;
  wire[5:0] T26;
  wire[25:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire T30;
  wire empty;
  wire T31;
  wire T32;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T33 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T34 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T35 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T19, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_payload_a_type, T17};
  assign T17 = {io_enq_bits_payload_union, io_enq_bits_payload_data};
  assign T18 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_is_builtin_type};
  assign T19 = {T21, T20};
  assign T20 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T21 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_union = T22;
  assign T22 = T11[8'h90:8'h80];
  assign io_deq_bits_payload_a_type = T23;
  assign T23 = T11[8'h93:8'h91];
  assign io_deq_bits_payload_is_builtin_type = T24;
  assign T24 = T11[8'h94];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h96:8'h95];
  assign io_deq_bits_payload_client_xact_id = T26;
  assign T26 = T11[8'h9c:8'h97];
  assign io_deq_bits_payload_addr_block = T27;
  assign T27 = T11[8'hb6:8'h9d];
  assign io_deq_bits_header_dst = T28;
  assign T28 = T11[8'hb9:8'hb7];
  assign io_deq_bits_header_src = T29;
  assign T29 = T11[8'hbc:8'hba];
  assign io_deq_valid = T30;
  assign T30 = empty ^ 1'h1;
  assign empty = ptr_match & T31;
  assign T31 = maybe_full ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_p_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T23;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T24;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[33:0] T11;
  reg [33:0] ram [1:0];
  wire[33:0] T12;
  wire[33:0] T13;
  wire[33:0] T14;
  wire[27:0] T15;
  wire[5:0] T16;
  wire[25:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_p_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_p_type};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T11[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T11[5'h1e:5'h1c];
  assign io_deq_bits_header_src = T19;
  assign T19 = T11[6'h21:5'h1f];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [5:0] io_enq_bits_payload_client_xact_id,
    input  io_enq_bits_payload_voluntary,
    input [2:0] io_enq_bits_payload_r_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[5:0] io_deq_bits_payload_client_xact_id,
    output io_deq_bits_payload_voluntary,
    output[2:0] io_deq_bits_payload_r_type,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[171:0] T11;
  reg [171:0] ram [1:0];
  wire[171:0] T12;
  wire[171:0] T13;
  wire[171:0] T14;
  wire[137:0] T15;
  wire[130:0] T16;
  wire[6:0] T17;
  wire[33:0] T18;
  wire[27:0] T19;
  wire[5:0] T20;
  wire[2:0] T21;
  wire T22;
  wire[5:0] T23;
  wire[25:0] T24;
  wire[1:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_r_type, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_voluntary};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T21;
  assign T21 = T11[8'h82:8'h80];
  assign io_deq_bits_payload_voluntary = T22;
  assign T22 = T11[8'h83];
  assign io_deq_bits_payload_client_xact_id = T23;
  assign T23 = T11[8'h89:8'h84];
  assign io_deq_bits_payload_addr_block = T24;
  assign T24 = T11[8'ha3:8'h8a];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'ha5:8'ha4];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'ha8:8'ha6];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'hab:8'ha9];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_16(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [5:0] io_enq_bits_payload_client_xact_id,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_enq_bits_payload_is_builtin_type,
    input [3:0] io_enq_bits_payload_g_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[5:0] io_deq_bits_payload_client_xact_id,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output io_deq_bits_payload_is_builtin_type,
    output[3:0] io_deq_bits_payload_g_type,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[150:0] T11;
  reg [150:0] ram [1:0];
  wire[150:0] T12;
  wire[150:0] T13;
  wire[150:0] T14;
  wire[136:0] T15;
  wire[131:0] T16;
  wire[4:0] T17;
  wire[13:0] T18;
  wire[7:0] T19;
  wire[5:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[3:0] T23;
  wire[5:0] T24;
  wire[1:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_g_type, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_manager_xact_id, io_enq_bits_payload_is_builtin_type};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_g_type = T21;
  assign T21 = T11[8'h83:8'h80];
  assign io_deq_bits_payload_is_builtin_type = T22;
  assign T22 = T11[8'h84];
  assign io_deq_bits_payload_manager_xact_id = T23;
  assign T23 = T11[8'h88:8'h85];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[8'h8e:8'h89];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h90:8'h8f];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'h93:8'h91];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'h96:8'h94];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_17(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[9:0] T11;
  reg [9:0] ram [1:0];
  wire[9:0] T12;
  wire[9:0] T13;
  wire[9:0] T14;
  wire[6:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_manager_xact_id = T10;
  assign T10 = T11[2'h3:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_header_src, T15};
  assign T15 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T16;
  assign T16 = T11[3'h6:3'h4];
  assign io_deq_bits_header_src = T17;
  assign T17 = T11[4'h9:3'h7];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module TileLinkEnqueuer_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [2:0] io_client_acquire_bits_header_src,
    input [2:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [5:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[2:0] io_client_grant_bits_header_src,
    output[2:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[5:0] io_client_grant_bits_payload_client_xact_id,
    output[3:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [2:0] io_client_finish_bits_header_src,
    input [2:0] io_client_finish_bits_header_dst,
    input [3:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[2:0] io_client_probe_bits_header_src,
    output[2:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [2:0] io_client_release_bits_header_src,
    input [2:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [5:0] io_client_release_bits_payload_client_xact_id,
    input  io_client_release_bits_payload_voluntary,
    input [2:0] io_client_release_bits_payload_r_type,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[2:0] io_manager_acquire_bits_header_src,
    output[2:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[5:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [2:0] io_manager_grant_bits_header_src,
    input [2:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [5:0] io_manager_grant_bits_payload_client_xact_id,
    input [3:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[2:0] io_manager_finish_bits_header_src,
    output[2:0] io_manager_finish_bits_header_dst,
    output[3:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [2:0] io_manager_probe_bits_header_src,
    input [2:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[2:0] io_manager_release_bits_header_src,
    output[2:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[5:0] io_manager_release_bits_payload_client_xact_id,
    output io_manager_release_bits_payload_voluntary,
    output[2:0] io_manager_release_bits_payload_r_type,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[2:0] Queue_io_deq_bits_header_src;
  wire[2:0] Queue_io_deq_bits_header_dst;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[5:0] Queue_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire Queue_io_deq_bits_payload_is_builtin_type;
  wire[2:0] Queue_io_deq_bits_payload_a_type;
  wire[16:0] Queue_io_deq_bits_payload_union;
  wire[127:0] Queue_io_deq_bits_payload_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[2:0] Queue_1_io_deq_bits_header_src;
  wire[2:0] Queue_1_io_deq_bits_header_dst;
  wire[25:0] Queue_1_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_1_io_deq_bits_payload_p_type;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[2:0] Queue_2_io_deq_bits_header_src;
  wire[2:0] Queue_2_io_deq_bits_header_dst;
  wire[1:0] Queue_2_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_2_io_deq_bits_payload_addr_block;
  wire[5:0] Queue_2_io_deq_bits_payload_client_xact_id;
  wire Queue_2_io_deq_bits_payload_voluntary;
  wire[2:0] Queue_2_io_deq_bits_payload_r_type;
  wire[127:0] Queue_2_io_deq_bits_payload_data;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[2:0] Queue_3_io_deq_bits_header_src;
  wire[2:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_payload_addr_beat;
  wire[5:0] Queue_3_io_deq_bits_payload_client_xact_id;
  wire[3:0] Queue_3_io_deq_bits_payload_manager_xact_id;
  wire Queue_3_io_deq_bits_payload_is_builtin_type;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire[127:0] Queue_3_io_deq_bits_payload_data;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[2:0] Queue_4_io_deq_bits_header_src;
  wire[2:0] Queue_4_io_deq_bits_header_dst;
  wire[3:0] Queue_4_io_deq_bits_payload_manager_xact_id;


  assign io_manager_release_bits_payload_data = Queue_2_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_r_type = Queue_2_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_voluntary = Queue_2_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_2_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_2_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_2_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_2_io_deq_valid;
  assign io_manager_probe_ready = Queue_1_io_enq_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = Queue_4_io_deq_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_finish_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_finish_valid = Queue_4_io_deq_valid;
  assign io_manager_grant_ready = Queue_3_io_enq_ready;
  assign io_manager_acquire_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = Queue_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = Queue_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_acquire_valid = Queue_io_deq_valid;
  assign io_client_release_ready = Queue_2_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = Queue_1_io_deq_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = Queue_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = Queue_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_header_src = Queue_1_io_deq_bits_header_src;
  assign io_client_probe_valid = Queue_1_io_deq_valid;
  assign io_client_finish_ready = Queue_4_io_enq_ready;
  assign io_client_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_client_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_client_grant_valid = Queue_3_io_deq_valid;
  assign io_client_acquire_ready = Queue_io_enq_ready;
  Queue_13 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_acquire_valid ),
       .io_enq_bits_header_src( io_client_acquire_bits_header_src ),
       .io_enq_bits_header_dst( io_client_acquire_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_acquire_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_acquire_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_acquire_bits_payload_addr_beat ),
       .io_enq_bits_payload_is_builtin_type( io_client_acquire_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_a_type( io_client_acquire_bits_payload_a_type ),
       .io_enq_bits_payload_union( io_client_acquire_bits_payload_union ),
       .io_enq_bits_payload_data( io_client_acquire_bits_payload_data ),
       .io_deq_ready( io_manager_acquire_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_is_builtin_type( Queue_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_a_type( Queue_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_union( Queue_io_deq_bits_payload_union ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_14 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( io_manager_probe_valid ),
       .io_enq_bits_header_src( io_manager_probe_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_probe_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_manager_probe_bits_payload_addr_block ),
       .io_enq_bits_payload_p_type( io_manager_probe_bits_payload_p_type ),
       .io_deq_ready( io_client_probe_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_1_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_p_type( Queue_1_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
  Queue_15 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_2_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_2_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_2_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_voluntary( Queue_2_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_r_type( Queue_2_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_data( Queue_2_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_16 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( io_manager_grant_valid ),
       .io_enq_bits_header_src( io_manager_grant_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_grant_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_manager_grant_bits_payload_addr_beat ),
       .io_enq_bits_payload_client_xact_id( io_manager_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( io_manager_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_is_builtin_type( io_manager_grant_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_g_type( io_manager_grant_bits_payload_g_type ),
       .io_enq_bits_payload_data( io_manager_grant_bits_payload_data ),
       .io_deq_ready( io_client_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_3_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_3_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_is_builtin_type( Queue_3_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_17 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( io_client_finish_valid ),
       .io_enq_bits_header_src( io_client_finish_bits_header_src ),
       .io_enq_bits_header_dst( io_client_finish_bits_header_dst ),
       .io_enq_bits_payload_manager_xact_id( io_client_finish_bits_payload_manager_xact_id ),
       .io_deq_ready( io_manager_finish_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_4_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
endmodule

module FinishUnit_1(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [2:0] io_grant_bits_header_src,
    input [2:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [5:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[5:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[2:0] io_finish_bits_header_src,
    output[2:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[2:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 3'h1;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [5:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[5:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [5:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[2:0] io_network_acquire_bits_header_src,
    output[2:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[5:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [2:0] io_network_grant_bits_header_src,
    input [2:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [5:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[2:0] io_network_finish_bits_header_src,
    output[2:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [2:0] io_network_probe_bits_header_src,
    input [2:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[2:0] io_network_release_bits_header_src,
    output[2:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[5:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[5:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[2:0] rel_with_header_bits_header_dst;
  wire[2:0] T8;
  wire T0;
  wire T1;
  wire[25:0] T2;
  wire[2:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[5:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[2:0] acq_with_header_bits_header_dst;
  wire[2:0] T9;
  wire T3;
  wire T4;
  wire[25:0] T5;
  wire[2:0] acq_with_header_bits_header_src;
  wire T6;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T7;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[5:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[2:0] finisher_io_finish_bits_header_src;
  wire[2:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = T8;
  assign T8 = {2'h0, T0};
  assign T0 = T1 == 1'h0;
  assign T1 = T2 < 26'h1000000;
  assign T2 = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 3'h1;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = T9;
  assign T9 = {2'h0, T3};
  assign T3 = T4 == 1'h0;
  assign T4 = T5 < 26'h1000000;
  assign T5 = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 3'h1;
  assign io_network_acquire_valid = T6;
  assign T6 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T7;
  assign T7 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_1 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module FinishUnit_2(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [2:0] io_grant_bits_header_src,
    input [2:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [5:0] io_grant_bits_payload_client_xact_id,
    input [3:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[5:0] io_refill_bits_client_xact_id,
    output[3:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[2:0] io_finish_bits_header_src,
    output[2:0] io_finish_bits_header_dst,
    output[3:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[3:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[3:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[2:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 3'h2;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_2(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [5:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[5:0] io_client_grant_bits_client_xact_id,
    output[3:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [5:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[2:0] io_network_acquire_bits_header_src,
    output[2:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[5:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [2:0] io_network_grant_bits_header_src,
    input [2:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [5:0] io_network_grant_bits_payload_client_xact_id,
    input [3:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[2:0] io_network_finish_bits_header_src,
    output[2:0] io_network_finish_bits_header_dst,
    output[3:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [2:0] io_network_probe_bits_header_src,
    input [2:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[2:0] io_network_release_bits_header_src,
    output[2:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[5:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[5:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[2:0] rel_with_header_bits_header_dst;
  wire[2:0] T8;
  wire T0;
  wire T1;
  wire[25:0] T2;
  wire[2:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[5:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[2:0] acq_with_header_bits_header_dst;
  wire[2:0] T9;
  wire T3;
  wire T4;
  wire[25:0] T5;
  wire[2:0] acq_with_header_bits_header_src;
  wire T6;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T7;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[5:0] finisher_io_refill_bits_client_xact_id;
  wire[3:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[2:0] finisher_io_finish_bits_header_src;
  wire[2:0] finisher_io_finish_bits_header_dst;
  wire[3:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = T8;
  assign T8 = {2'h0, T0};
  assign T0 = T1 == 1'h0;
  assign T1 = T2 < 26'h1000000;
  assign T2 = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 3'h2;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = T9;
  assign T9 = {2'h0, T3};
  assign T3 = T4 == 1'h0;
  assign T4 = T5 < 26'h1000000;
  assign T5 = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 3'h2;
  assign io_network_acquire_valid = T6;
  assign T6 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T7;
  assign T7 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_2 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module ManagerTileLinkNetworkPort_0(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output[5:0] io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output[127:0] io_manager_acquire_bits_data,
    output[1:0] io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [5:0] io_manager_grant_bits_client_xact_id,
    input [3:0] io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input [127:0] io_manager_grant_bits_data,
    input [1:0] io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[3:0] io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input [1:0] io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_addr_beat,
    output[25:0] io_manager_release_bits_addr_block,
    output[5:0] io_manager_release_bits_client_xact_id,
    output io_manager_release_bits_voluntary,
    output[2:0] io_manager_release_bits_r_type,
    output[127:0] io_manager_release_bits_data,
    output[1:0] io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input [2:0] io_network_acquire_bits_header_src,
    input [2:0] io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input [5:0] io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output[2:0] io_network_grant_bits_header_src,
    output[2:0] io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[5:0] io_network_grant_bits_payload_client_xact_id,
    output[3:0] io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output[127:0] io_network_grant_bits_payload_data,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input [2:0] io_network_finish_bits_header_src,
    input [2:0] io_network_finish_bits_header_dst,
    input [3:0] io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output[2:0] io_network_probe_bits_header_src,
    output[2:0] io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input [2:0] io_network_release_bits_header_src,
    input [2:0] io_network_release_bits_header_dst,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [25:0] io_network_release_bits_payload_addr_block,
    input [5:0] io_network_release_bits_payload_client_xact_id,
    input  io_network_release_bits_payload_voluntary,
    input [2:0] io_network_release_bits_payload_r_type,
    input [127:0] io_network_release_bits_payload_data
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire[2:0] T3;
  wire[2:0] T36;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[127:0] T7;
  wire[3:0] T8;
  wire T9;
  wire[3:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire[2:0] T13;
  wire[2:0] T37;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire[1:0] T38;
  wire[127:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[5:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T39;
  wire[127:0] T28;
  wire[16:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[5:0] T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = T36;
  assign T36 = {1'h0, io_manager_probe_bits_client_id};
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 3'h0;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_data = T7;
  assign T7 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_g_type = T8;
  assign T8 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T9;
  assign T9 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T10;
  assign T10 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T11;
  assign T11 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = T37;
  assign T37 = {1'h0, io_manager_grant_bits_client_id};
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 3'h0;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = T38;
  assign T38 = io_network_release_bits_header_src[1'h1:1'h0];
  assign io_manager_release_bits_data = T17;
  assign T17 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_r_type = T18;
  assign T18 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_voluntary = T19;
  assign T19 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_client_xact_id = T20;
  assign T20 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T21;
  assign T21 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_bits_addr_beat = T22;
  assign T22 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = T39;
  assign T39 = io_network_acquire_bits_header_src[1'h1:1'h0];
  assign io_manager_acquire_bits_data = T28;
  assign T28 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_union = T29;
  assign T29 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T30;
  assign T30 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T31;
  assign T31 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module Queue_18(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_header_src,
    input [2:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [5:0] io_enq_bits_payload_client_xact_id,
    input  io_enq_bits_payload_voluntary,
    input [2:0] io_enq_bits_payload_r_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_header_src,
    output[2:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[5:0] io_deq_bits_payload_client_xact_id,
    output io_deq_bits_payload_voluntary,
    output[2:0] io_deq_bits_payload_r_type,
    output[127:0] io_deq_bits_payload_data,
    output io_count
);

  wire T23;
  wire[1:0] T0;
  reg  full;
  wire T24;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[171:0] T4;
  reg [171:0] ram [0:0];
  wire[171:0] T5;
  wire[171:0] T6;
  wire[171:0] T7;
  wire[137:0] T8;
  wire[130:0] T9;
  wire[6:0] T10;
  wire[33:0] T11;
  wire[27:0] T12;
  wire[5:0] T13;
  wire[2:0] T14;
  wire T15;
  wire[5:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire empty;
  wire T22;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T23;
  assign T23 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T24 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_payload_r_type, io_enq_bits_payload_data};
  assign T10 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_voluntary};
  assign T11 = {T13, T12};
  assign T12 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T13 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T14;
  assign T14 = T4[8'h82:8'h80];
  assign io_deq_bits_payload_voluntary = T15;
  assign T15 = T4[8'h83];
  assign io_deq_bits_payload_client_xact_id = T16;
  assign T16 = T4[8'h89:8'h84];
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T4[8'ha3:8'h8a];
  assign io_deq_bits_payload_addr_beat = T18;
  assign T18 = T4[8'ha5:8'ha4];
  assign io_deq_bits_header_dst = T19;
  assign T19 = T4[8'ha8:8'ha6];
  assign io_deq_bits_header_src = T20;
  assign T20 = T4[8'hab:8'ha9];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module TileLinkEnqueuer_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [2:0] io_client_acquire_bits_header_src,
    input [2:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [5:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[2:0] io_client_grant_bits_header_src,
    output[2:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[5:0] io_client_grant_bits_payload_client_xact_id,
    output[3:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [2:0] io_client_finish_bits_header_src,
    input [2:0] io_client_finish_bits_header_dst,
    input [3:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[2:0] io_client_probe_bits_header_src,
    output[2:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [2:0] io_client_release_bits_header_src,
    input [2:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [5:0] io_client_release_bits_payload_client_xact_id,
    input  io_client_release_bits_payload_voluntary,
    input [2:0] io_client_release_bits_payload_r_type,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[2:0] io_manager_acquire_bits_header_src,
    output[2:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[5:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [2:0] io_manager_grant_bits_header_src,
    input [2:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [5:0] io_manager_grant_bits_payload_client_xact_id,
    input [3:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[2:0] io_manager_finish_bits_header_src,
    output[2:0] io_manager_finish_bits_header_dst,
    output[3:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [2:0] io_manager_probe_bits_header_src,
    input [2:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[2:0] io_manager_release_bits_header_src,
    output[2:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[5:0] io_manager_release_bits_payload_client_xact_id,
    output io_manager_release_bits_payload_voluntary,
    output[2:0] io_manager_release_bits_payload_r_type,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[2:0] Queue_io_deq_bits_header_src;
  wire[2:0] Queue_io_deq_bits_header_dst;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[5:0] Queue_io_deq_bits_payload_client_xact_id;
  wire Queue_io_deq_bits_payload_voluntary;
  wire[2:0] Queue_io_deq_bits_payload_r_type;
  wire[127:0] Queue_io_deq_bits_payload_data;


  assign io_manager_release_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_r_type = Queue_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_voluntary = Queue_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_io_deq_valid;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_client_release_ready = Queue_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_acquire_ready = io_manager_acquire_ready;
  Queue_18 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_voluntary( Queue_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_r_type( Queue_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
endmodule

module ManagerTileLinkNetworkPort_1(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output[5:0] io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output[127:0] io_manager_acquire_bits_data,
    output[1:0] io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [5:0] io_manager_grant_bits_client_xact_id,
    input [3:0] io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input [127:0] io_manager_grant_bits_data,
    input [1:0] io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[3:0] io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input [1:0] io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_addr_beat,
    output[25:0] io_manager_release_bits_addr_block,
    output[5:0] io_manager_release_bits_client_xact_id,
    output io_manager_release_bits_voluntary,
    output[2:0] io_manager_release_bits_r_type,
    output[127:0] io_manager_release_bits_data,
    output[1:0] io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input [2:0] io_network_acquire_bits_header_src,
    input [2:0] io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input [5:0] io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output[2:0] io_network_grant_bits_header_src,
    output[2:0] io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[5:0] io_network_grant_bits_payload_client_xact_id,
    output[3:0] io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output[127:0] io_network_grant_bits_payload_data,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input [2:0] io_network_finish_bits_header_src,
    input [2:0] io_network_finish_bits_header_dst,
    input [3:0] io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output[2:0] io_network_probe_bits_header_src,
    output[2:0] io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input [2:0] io_network_release_bits_header_src,
    input [2:0] io_network_release_bits_header_dst,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [25:0] io_network_release_bits_payload_addr_block,
    input [5:0] io_network_release_bits_payload_client_xact_id,
    input  io_network_release_bits_payload_voluntary,
    input [2:0] io_network_release_bits_payload_r_type,
    input [127:0] io_network_release_bits_payload_data
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire[2:0] T3;
  wire[2:0] T36;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire[127:0] T7;
  wire[3:0] T8;
  wire T9;
  wire[3:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire[2:0] T13;
  wire[2:0] T37;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire[1:0] T38;
  wire[127:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[5:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T39;
  wire[127:0] T28;
  wire[16:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[5:0] T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = T36;
  assign T36 = {1'h0, io_manager_probe_bits_client_id};
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 3'h1;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_data = T7;
  assign T7 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_g_type = T8;
  assign T8 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T9;
  assign T9 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T10;
  assign T10 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T11;
  assign T11 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = T37;
  assign T37 = {1'h0, io_manager_grant_bits_client_id};
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 3'h1;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = T38;
  assign T38 = io_network_release_bits_header_src[1'h1:1'h0];
  assign io_manager_release_bits_data = T17;
  assign T17 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_r_type = T18;
  assign T18 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_voluntary = T19;
  assign T19 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_client_xact_id = T20;
  assign T20 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T21;
  assign T21 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_bits_addr_beat = T22;
  assign T22 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = T39;
  assign T39 = io_network_acquire_bits_header_src[1'h1:1'h0];
  assign io_manager_acquire_bits_data = T28;
  assign T28 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_union = T29;
  assign T29 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T30;
  assign T30 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T31;
  assign T31 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module LockingRRArbiter_5(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input  io_in_4_bits_payload_is_builtin_type,
    input [2:0] io_in_4_bits_payload_a_type,
    input [16:0] io_in_4_bits_payload_union,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input  io_in_3_bits_payload_is_builtin_type,
    input [2:0] io_in_3_bits_payload_a_type,
    input [16:0] io_in_3_bits_payload_union,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input  io_in_2_bits_payload_is_builtin_type,
    input [2:0] io_in_2_bits_payload_a_type,
    input [16:0] io_in_2_bits_payload_union,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input  io_in_1_bits_payload_is_builtin_type,
    input [2:0] io_in_1_bits_payload_a_type,
    input [16:0] io_in_1_bits_payload_union,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input  io_in_0_bits_payload_is_builtin_type,
    input [2:0] io_in_0_bits_payload_a_type,
    input [16:0] io_in_0_bits_payload_union,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_header_src,
    output[2:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output[5:0] io_out_bits_payload_client_xact_id,
    output[1:0] io_out_bits_payload_addr_beat,
    output io_out_bits_payload_is_builtin_type,
    output[2:0] io_out_bits_payload_a_type,
    output[16:0] io_out_bits_payload_union,
    output[127:0] io_out_bits_payload_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T207;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T208;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  locked;
  wire T209;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  reg [1:0] R38;
  wire[1:0] T210;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire[127:0] T42;
  wire[127:0] T43;
  wire[127:0] T44;
  wire T45;
  wire[2:0] T46;
  wire[127:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[16:0] T51;
  wire[16:0] T52;
  wire[16:0] T53;
  wire T54;
  wire[16:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[2:0] T60;
  wire[2:0] T61;
  wire T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire T78;
  wire[1:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire[5:0] T83;
  wire[5:0] T84;
  wire[5:0] T85;
  wire T86;
  wire[5:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[25:0] T91;
  wire[25:0] T92;
  wire[25:0] T93;
  wire T94;
  wire[25:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[2:0] T99;
  wire[2:0] T100;
  wire[2:0] T101;
  wire T102;
  wire[2:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire T110;
  wire[2:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R38 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T207 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T208 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T32 & T30;
  assign T30 = io_out_bits_payload_is_builtin_type & T31;
  assign T31 = 3'h3 == io_out_bits_payload_a_type;
  assign T32 = io_out_valid & io_out_ready;
  assign T209 = reset ? 1'h0 : T33;
  assign T33 = T40 ? 1'h0 : T34;
  assign T34 = T29 ? T35 : locked;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 == 2'h0;
  assign T37 = R38 + 2'h1;
  assign T210 = reset ? 2'h0 : T39;
  assign T39 = T29 ? T37 : R38;
  assign T40 = T32 & T41;
  assign T41 = T30 ^ 1'h1;
  assign io_out_bits_payload_data = T42;
  assign T42 = T50 ? io_in_4_bits_payload_data : T43;
  assign T43 = T49 ? T47 : T44;
  assign T44 = T45 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T45 = T46[1'h0];
  assign T46 = chosen;
  assign T47 = T48 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T48 = T46[1'h0];
  assign T49 = T46[1'h1];
  assign T50 = T46[2'h2];
  assign io_out_bits_payload_union = T51;
  assign T51 = T58 ? io_in_4_bits_payload_union : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign T54 = T46[1'h0];
  assign T55 = T56 ? io_in_3_bits_payload_union : io_in_2_bits_payload_union;
  assign T56 = T46[1'h0];
  assign T57 = T46[1'h1];
  assign T58 = T46[2'h2];
  assign io_out_bits_payload_a_type = T59;
  assign T59 = T66 ? io_in_4_bits_payload_a_type : T60;
  assign T60 = T65 ? T63 : T61;
  assign T61 = T62 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T62 = T46[1'h0];
  assign T63 = T64 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T64 = T46[1'h0];
  assign T65 = T46[1'h1];
  assign T66 = T46[2'h2];
  assign io_out_bits_payload_is_builtin_type = T67;
  assign T67 = T74 ? io_in_4_bits_payload_is_builtin_type : T68;
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign T70 = T46[1'h0];
  assign T71 = T72 ? io_in_3_bits_payload_is_builtin_type : io_in_2_bits_payload_is_builtin_type;
  assign T72 = T46[1'h0];
  assign T73 = T46[1'h1];
  assign T74 = T46[2'h2];
  assign io_out_bits_payload_addr_beat = T75;
  assign T75 = T82 ? io_in_4_bits_payload_addr_beat : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T78 = T46[1'h0];
  assign T79 = T80 ? io_in_3_bits_payload_addr_beat : io_in_2_bits_payload_addr_beat;
  assign T80 = T46[1'h0];
  assign T81 = T46[1'h1];
  assign T82 = T46[2'h2];
  assign io_out_bits_payload_client_xact_id = T83;
  assign T83 = T90 ? io_in_4_bits_payload_client_xact_id : T84;
  assign T84 = T89 ? T87 : T85;
  assign T85 = T86 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T86 = T46[1'h0];
  assign T87 = T88 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T88 = T46[1'h0];
  assign T89 = T46[1'h1];
  assign T90 = T46[2'h2];
  assign io_out_bits_payload_addr_block = T91;
  assign T91 = T98 ? io_in_4_bits_payload_addr_block : T92;
  assign T92 = T97 ? T95 : T93;
  assign T93 = T94 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T94 = T46[1'h0];
  assign T95 = T96 ? io_in_3_bits_payload_addr_block : io_in_2_bits_payload_addr_block;
  assign T96 = T46[1'h0];
  assign T97 = T46[1'h1];
  assign T98 = T46[2'h2];
  assign io_out_bits_header_dst = T99;
  assign T99 = T106 ? io_in_4_bits_header_dst : T100;
  assign T100 = T105 ? T103 : T101;
  assign T101 = T102 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T102 = T46[1'h0];
  assign T103 = T104 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T104 = T46[1'h0];
  assign T105 = T46[1'h1];
  assign T106 = T46[2'h2];
  assign io_out_bits_header_src = T107;
  assign T107 = T114 ? io_in_4_bits_header_src : T108;
  assign T108 = T113 ? T111 : T109;
  assign T109 = T110 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T110 = T46[1'h0];
  assign T111 = T112 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T112 = T46[1'h0];
  assign T113 = T46[1'h1];
  assign T114 = T46[2'h2];
  assign io_out_valid = T115;
  assign T115 = T122 ? io_in_4_valid : T116;
  assign T116 = T121 ? T119 : T117;
  assign T117 = T118 ? io_in_1_valid : io_in_0_valid;
  assign T118 = T46[1'h0];
  assign T119 = T120 ? io_in_3_valid : io_in_2_valid;
  assign T120 = T46[1'h0];
  assign T121 = T46[1'h1];
  assign T122 = T46[2'h2];
  assign io_in_0_ready = T123;
  assign T123 = T124 & io_out_ready;
  assign T124 = locked ? T142 : T125;
  assign T125 = T141 | T126;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T130 | T128;
  assign T128 = io_in_4_valid & T129;
  assign T129 = last_grant < 3'h4;
  assign T130 = T133 | T131;
  assign T131 = io_in_3_valid & T132;
  assign T132 = last_grant < 3'h3;
  assign T133 = T136 | T134;
  assign T134 = io_in_2_valid & T135;
  assign T135 = last_grant < 3'h2;
  assign T136 = T139 | T137;
  assign T137 = io_in_1_valid & T138;
  assign T138 = last_grant < 3'h1;
  assign T139 = io_in_0_valid & T140;
  assign T140 = last_grant < 3'h0;
  assign T141 = last_grant < 3'h0;
  assign T142 = lockIdx == 3'h0;
  assign io_in_1_ready = T143;
  assign T143 = T144 & io_out_ready;
  assign T144 = locked ? T155 : T145;
  assign T145 = T152 | T146;
  assign T146 = T147 ^ 1'h1;
  assign T147 = T148 | io_in_0_valid;
  assign T148 = T149 | T128;
  assign T149 = T150 | T131;
  assign T150 = T151 | T134;
  assign T151 = T139 | T137;
  assign T152 = T154 & T153;
  assign T153 = last_grant < 3'h1;
  assign T154 = T139 ^ 1'h1;
  assign T155 = lockIdx == 3'h1;
  assign io_in_2_ready = T156;
  assign T156 = T157 & io_out_ready;
  assign T157 = locked ? T170 : T158;
  assign T158 = T166 | T159;
  assign T159 = T160 ^ 1'h1;
  assign T160 = T161 | io_in_1_valid;
  assign T161 = T162 | io_in_0_valid;
  assign T162 = T163 | T128;
  assign T163 = T164 | T131;
  assign T164 = T165 | T134;
  assign T165 = T139 | T137;
  assign T166 = T168 & T167;
  assign T167 = last_grant < 3'h2;
  assign T168 = T169 ^ 1'h1;
  assign T169 = T139 | T137;
  assign T170 = lockIdx == 3'h2;
  assign io_in_3_ready = T171;
  assign T171 = T172 & io_out_ready;
  assign T172 = locked ? T187 : T173;
  assign T173 = T182 | T174;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T176 | io_in_2_valid;
  assign T176 = T177 | io_in_1_valid;
  assign T177 = T178 | io_in_0_valid;
  assign T178 = T179 | T128;
  assign T179 = T180 | T131;
  assign T180 = T181 | T134;
  assign T181 = T139 | T137;
  assign T182 = T184 & T183;
  assign T183 = last_grant < 3'h3;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T186 | T134;
  assign T186 = T139 | T137;
  assign T187 = lockIdx == 3'h3;
  assign io_in_4_ready = T188;
  assign T188 = T189 & io_out_ready;
  assign T189 = locked ? T206 : T190;
  assign T190 = T200 | T191;
  assign T191 = T192 ^ 1'h1;
  assign T192 = T193 | io_in_3_valid;
  assign T193 = T194 | io_in_2_valid;
  assign T194 = T195 | io_in_1_valid;
  assign T195 = T196 | io_in_0_valid;
  assign T196 = T197 | T128;
  assign T197 = T198 | T131;
  assign T198 = T199 | T134;
  assign T199 = T139 | T137;
  assign T200 = T202 & T201;
  assign T201 = last_grant < 3'h4;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T204 | T131;
  assign T204 = T205 | T134;
  assign T205 = T139 | T137;
  assign T206 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T40) begin
      locked <= 1'h0;
    end else if(T29) begin
      locked <= T35;
    end
    if(reset) begin
      R38 <= 2'h0;
    end else if(T29) begin
      R38 <= T37;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input  io_in_4_bits_payload_is_builtin_type,
    input [2:0] io_in_4_bits_payload_a_type,
    input [16:0] io_in_4_bits_payload_union,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input  io_in_3_bits_payload_is_builtin_type,
    input [2:0] io_in_3_bits_payload_a_type,
    input [16:0] io_in_3_bits_payload_union,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input  io_in_2_bits_payload_is_builtin_type,
    input [2:0] io_in_2_bits_payload_a_type,
    input [16:0] io_in_2_bits_payload_union,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input  io_in_1_bits_payload_is_builtin_type,
    input [2:0] io_in_1_bits_payload_a_type,
    input [16:0] io_in_1_bits_payload_union,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input  io_in_0_bits_payload_is_builtin_type,
    input [2:0] io_in_0_bits_payload_a_type,
    input [16:0] io_in_0_bits_payload_union,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_4_ready,
    output io_out_4_valid,
    output[2:0] io_out_4_bits_header_src,
    output[2:0] io_out_4_bits_header_dst,
    output[25:0] io_out_4_bits_payload_addr_block,
    output[5:0] io_out_4_bits_payload_client_xact_id,
    output[1:0] io_out_4_bits_payload_addr_beat,
    output io_out_4_bits_payload_is_builtin_type,
    output[2:0] io_out_4_bits_payload_a_type,
    output[16:0] io_out_4_bits_payload_union,
    output[127:0] io_out_4_bits_payload_data,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[2:0] io_out_3_bits_header_src,
    output[2:0] io_out_3_bits_header_dst,
    output[25:0] io_out_3_bits_payload_addr_block,
    output[5:0] io_out_3_bits_payload_client_xact_id,
    output[1:0] io_out_3_bits_payload_addr_beat,
    output io_out_3_bits_payload_is_builtin_type,
    output[2:0] io_out_3_bits_payload_a_type,
    output[16:0] io_out_3_bits_payload_union,
    output[127:0] io_out_3_bits_payload_data,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[2:0] io_out_2_bits_header_src,
    output[2:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr_block,
    output[5:0] io_out_2_bits_payload_client_xact_id,
    output[1:0] io_out_2_bits_payload_addr_beat,
    output io_out_2_bits_payload_is_builtin_type,
    output[2:0] io_out_2_bits_payload_a_type,
    output[16:0] io_out_2_bits_payload_union,
    output[127:0] io_out_2_bits_payload_data,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[2:0] io_out_1_bits_header_src,
    output[2:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr_block,
    output[5:0] io_out_1_bits_payload_client_xact_id,
    output[1:0] io_out_1_bits_payload_addr_beat,
    output io_out_1_bits_payload_is_builtin_type,
    output[2:0] io_out_1_bits_payload_a_type,
    output[16:0] io_out_1_bits_payload_union,
    output[127:0] io_out_1_bits_payload_data,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[2:0] io_out_0_bits_header_src,
    output[2:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr_block,
    output[5:0] io_out_0_bits_payload_client_xact_id,
    output[1:0] io_out_0_bits_payload_addr_beat,
    output io_out_0_bits_payload_is_builtin_type,
    output[2:0] io_out_0_bits_payload_a_type,
    output[16:0] io_out_0_bits_payload_union,
    output[127:0] io_out_0_bits_payload_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[2:0] LockingRRArbiter_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_1_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_1_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire LockingRRArbiter_2_io_in_4_ready;
  wire LockingRRArbiter_2_io_in_3_ready;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_2_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_2_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire LockingRRArbiter_3_io_in_4_ready;
  wire LockingRRArbiter_3_io_in_3_ready;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_3_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_3_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire LockingRRArbiter_4_io_in_4_ready;
  wire LockingRRArbiter_4_io_in_3_ready;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_4_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_4_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_4_io_out_bits_payload_data;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 3'h4;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 3'h4;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 3'h4;
  assign T6 = io_in_3_valid & T7;
  assign T7 = io_in_3_bits_header_dst == 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = io_in_4_bits_header_dst == 3'h4;
  assign T10 = io_in_0_valid & T11;
  assign T11 = io_in_0_bits_header_dst == 3'h3;
  assign T12 = io_in_1_valid & T13;
  assign T13 = io_in_1_bits_header_dst == 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = io_in_2_bits_header_dst == 3'h3;
  assign T16 = io_in_3_valid & T17;
  assign T17 = io_in_3_bits_header_dst == 3'h3;
  assign T18 = io_in_4_valid & T19;
  assign T19 = io_in_4_bits_header_dst == 3'h3;
  assign T20 = io_in_0_valid & T21;
  assign T21 = io_in_0_bits_header_dst == 3'h2;
  assign T22 = io_in_1_valid & T23;
  assign T23 = io_in_1_bits_header_dst == 3'h2;
  assign T24 = io_in_2_valid & T25;
  assign T25 = io_in_2_bits_header_dst == 3'h2;
  assign T26 = io_in_3_valid & T27;
  assign T27 = io_in_3_bits_header_dst == 3'h2;
  assign T28 = io_in_4_valid & T29;
  assign T29 = io_in_4_bits_header_dst == 3'h2;
  assign T30 = io_in_0_valid & T31;
  assign T31 = io_in_0_bits_header_dst == 3'h1;
  assign T32 = io_in_1_valid & T33;
  assign T33 = io_in_1_bits_header_dst == 3'h1;
  assign T34 = io_in_2_valid & T35;
  assign T35 = io_in_2_bits_header_dst == 3'h1;
  assign T36 = io_in_3_valid & T37;
  assign T37 = io_in_3_bits_header_dst == 3'h1;
  assign T38 = io_in_4_valid & T39;
  assign T39 = io_in_4_bits_header_dst == 3'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = io_in_0_bits_header_dst == 3'h0;
  assign T42 = io_in_1_valid & T43;
  assign T43 = io_in_1_bits_header_dst == 3'h0;
  assign T44 = io_in_2_valid & T45;
  assign T45 = io_in_2_bits_header_dst == 3'h0;
  assign T46 = io_in_3_valid & T47;
  assign T47 = io_in_3_bits_header_dst == 3'h0;
  assign T48 = io_in_4_valid & T49;
  assign T49 = io_in_4_bits_header_dst == 3'h0;
  assign io_out_0_bits_payload_data = LockingRRArbiter_io_out_bits_payload_data;
  assign io_out_0_bits_payload_union = LockingRRArbiter_io_out_bits_payload_union;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_is_builtin_type = LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_addr_beat = LockingRRArbiter_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_block = LockingRRArbiter_io_out_bits_payload_addr_block;
  assign io_out_0_bits_header_dst = LockingRRArbiter_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_io_out_valid;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_union = LockingRRArbiter_1_io_out_bits_payload_union;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_is_builtin_type = LockingRRArbiter_1_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_addr_beat = LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_block = LockingRRArbiter_1_io_out_bits_payload_addr_block;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_union = LockingRRArbiter_2_io_out_bits_payload_union;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_is_builtin_type = LockingRRArbiter_2_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_addr_beat = LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_block = LockingRRArbiter_2_io_out_bits_payload_addr_block;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_out_3_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_3_bits_payload_union = LockingRRArbiter_3_io_out_bits_payload_union;
  assign io_out_3_bits_payload_a_type = LockingRRArbiter_3_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_is_builtin_type = LockingRRArbiter_3_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_addr_beat = LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_block = LockingRRArbiter_3_io_out_bits_payload_addr_block;
  assign io_out_3_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_3_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_3_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_4_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_4_bits_payload_union = LockingRRArbiter_4_io_out_bits_payload_union;
  assign io_out_4_bits_payload_a_type = LockingRRArbiter_4_io_out_bits_payload_a_type;
  assign io_out_4_bits_payload_is_builtin_type = LockingRRArbiter_4_io_out_bits_payload_is_builtin_type;
  assign io_out_4_bits_payload_addr_beat = LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_addr_block = LockingRRArbiter_4_io_out_bits_payload_addr_block;
  assign io_out_4_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_4_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_4_valid = LockingRRArbiter_4_io_out_valid;
  assign io_in_0_ready = T50;
  assign T50 = T54 | T51;
  assign T51 = T52;
  assign T52 = LockingRRArbiter_4_io_in_0_ready & T53;
  assign T53 = io_in_0_bits_header_dst == 3'h4;
  assign T54 = T58 | T55;
  assign T55 = T56;
  assign T56 = LockingRRArbiter_3_io_in_0_ready & T57;
  assign T57 = io_in_0_bits_header_dst == 3'h3;
  assign T58 = T62 | T59;
  assign T59 = T60;
  assign T60 = LockingRRArbiter_2_io_in_0_ready & T61;
  assign T61 = io_in_0_bits_header_dst == 3'h2;
  assign T62 = T66 | T63;
  assign T63 = T64;
  assign T64 = LockingRRArbiter_1_io_in_0_ready & T65;
  assign T65 = io_in_0_bits_header_dst == 3'h1;
  assign T66 = T67;
  assign T67 = LockingRRArbiter_io_in_0_ready & T68;
  assign T68 = io_in_0_bits_header_dst == 3'h0;
  assign io_in_1_ready = T69;
  assign T69 = T73 | T70;
  assign T70 = T71;
  assign T71 = LockingRRArbiter_4_io_in_1_ready & T72;
  assign T72 = io_in_1_bits_header_dst == 3'h4;
  assign T73 = T77 | T74;
  assign T74 = T75;
  assign T75 = LockingRRArbiter_3_io_in_1_ready & T76;
  assign T76 = io_in_1_bits_header_dst == 3'h3;
  assign T77 = T81 | T78;
  assign T78 = T79;
  assign T79 = LockingRRArbiter_2_io_in_1_ready & T80;
  assign T80 = io_in_1_bits_header_dst == 3'h2;
  assign T81 = T85 | T82;
  assign T82 = T83;
  assign T83 = LockingRRArbiter_1_io_in_1_ready & T84;
  assign T84 = io_in_1_bits_header_dst == 3'h1;
  assign T85 = T86;
  assign T86 = LockingRRArbiter_io_in_1_ready & T87;
  assign T87 = io_in_1_bits_header_dst == 3'h0;
  assign io_in_2_ready = T88;
  assign T88 = T92 | T89;
  assign T89 = T90;
  assign T90 = LockingRRArbiter_4_io_in_2_ready & T91;
  assign T91 = io_in_2_bits_header_dst == 3'h4;
  assign T92 = T96 | T93;
  assign T93 = T94;
  assign T94 = LockingRRArbiter_3_io_in_2_ready & T95;
  assign T95 = io_in_2_bits_header_dst == 3'h3;
  assign T96 = T100 | T97;
  assign T97 = T98;
  assign T98 = LockingRRArbiter_2_io_in_2_ready & T99;
  assign T99 = io_in_2_bits_header_dst == 3'h2;
  assign T100 = T104 | T101;
  assign T101 = T102;
  assign T102 = LockingRRArbiter_1_io_in_2_ready & T103;
  assign T103 = io_in_2_bits_header_dst == 3'h1;
  assign T104 = T105;
  assign T105 = LockingRRArbiter_io_in_2_ready & T106;
  assign T106 = io_in_2_bits_header_dst == 3'h0;
  assign io_in_3_ready = T107;
  assign T107 = T111 | T108;
  assign T108 = T109;
  assign T109 = LockingRRArbiter_4_io_in_3_ready & T110;
  assign T110 = io_in_3_bits_header_dst == 3'h4;
  assign T111 = T115 | T112;
  assign T112 = T113;
  assign T113 = LockingRRArbiter_3_io_in_3_ready & T114;
  assign T114 = io_in_3_bits_header_dst == 3'h3;
  assign T115 = T119 | T116;
  assign T116 = T117;
  assign T117 = LockingRRArbiter_2_io_in_3_ready & T118;
  assign T118 = io_in_3_bits_header_dst == 3'h2;
  assign T119 = T123 | T120;
  assign T120 = T121;
  assign T121 = LockingRRArbiter_1_io_in_3_ready & T122;
  assign T122 = io_in_3_bits_header_dst == 3'h1;
  assign T123 = T124;
  assign T124 = LockingRRArbiter_io_in_3_ready & T125;
  assign T125 = io_in_3_bits_header_dst == 3'h0;
  assign io_in_4_ready = T126;
  assign T126 = T130 | T127;
  assign T127 = T128;
  assign T128 = LockingRRArbiter_4_io_in_4_ready & T129;
  assign T129 = io_in_4_bits_header_dst == 3'h4;
  assign T130 = T134 | T131;
  assign T131 = T132;
  assign T132 = LockingRRArbiter_3_io_in_4_ready & T133;
  assign T133 = io_in_4_bits_header_dst == 3'h3;
  assign T134 = T138 | T135;
  assign T135 = T136;
  assign T136 = LockingRRArbiter_2_io_in_4_ready & T137;
  assign T137 = io_in_4_bits_header_dst == 3'h2;
  assign T138 = T142 | T139;
  assign T139 = T140;
  assign T140 = LockingRRArbiter_1_io_in_4_ready & T141;
  assign T141 = io_in_4_bits_header_dst == 3'h1;
  assign T142 = T143;
  assign T143 = LockingRRArbiter_io_in_4_ready & T144;
  assign T144 = io_in_4_bits_header_dst == 3'h0;
  LockingRRArbiter_5 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( T48 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_a_type( io_in_4_bits_payload_a_type ),
       .io_in_4_bits_payload_union( io_in_4_bits_payload_union ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( T46 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_a_type( io_in_3_bits_payload_a_type ),
       .io_in_3_bits_payload_union( io_in_3_bits_payload_union ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( T44 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_union( io_in_2_bits_payload_union ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( T42 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_union( io_in_1_bits_payload_union ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_union( io_in_0_bits_payload_union ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_5 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( T38 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_a_type( io_in_4_bits_payload_a_type ),
       .io_in_4_bits_payload_union( io_in_4_bits_payload_union ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( T36 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_a_type( io_in_3_bits_payload_a_type ),
       .io_in_3_bits_payload_union( io_in_3_bits_payload_union ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T34 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_union( io_in_2_bits_payload_union ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T32 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_union( io_in_1_bits_payload_union ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T30 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_union( io_in_0_bits_payload_union ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_1_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_1_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_5 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( T28 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_a_type( io_in_4_bits_payload_a_type ),
       .io_in_4_bits_payload_union( io_in_4_bits_payload_union ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( T26 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_a_type( io_in_3_bits_payload_a_type ),
       .io_in_3_bits_payload_union( io_in_3_bits_payload_union ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T24 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_union( io_in_2_bits_payload_union ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T22 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_union( io_in_1_bits_payload_union ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_union( io_in_0_bits_payload_union ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_2_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_2_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_2_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_2_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_5 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( T18 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_a_type( io_in_4_bits_payload_a_type ),
       .io_in_4_bits_payload_union( io_in_4_bits_payload_union ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( T16 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_a_type( io_in_3_bits_payload_a_type ),
       .io_in_3_bits_payload_union( io_in_3_bits_payload_union ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T14 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_union( io_in_2_bits_payload_union ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T12 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_union( io_in_1_bits_payload_union ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T10 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_union( io_in_0_bits_payload_union ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_3_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_3_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_3_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_3_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_3_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_3_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_5 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_4_io_in_4_ready ),
       .io_in_4_valid( T8 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_a_type( io_in_4_bits_payload_a_type ),
       .io_in_4_bits_payload_union( io_in_4_bits_payload_union ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_4_io_in_3_ready ),
       .io_in_3_valid( T6 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_a_type( io_in_3_bits_payload_a_type ),
       .io_in_3_bits_payload_union( io_in_3_bits_payload_union ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_union( io_in_2_bits_payload_union ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_union( io_in_1_bits_payload_union ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_union( io_in_0_bits_payload_union ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_4_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_4_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_4_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_4_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_4_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_4_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_6(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input  io_in_4_bits_payload_voluntary,
    input [2:0] io_in_4_bits_payload_r_type,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input  io_in_3_bits_payload_voluntary,
    input [2:0] io_in_3_bits_payload_r_type,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input  io_in_2_bits_payload_voluntary,
    input [2:0] io_in_2_bits_payload_r_type,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input  io_in_1_bits_payload_voluntary,
    input [2:0] io_in_1_bits_payload_r_type,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input  io_in_0_bits_payload_voluntary,
    input [2:0] io_in_0_bits_payload_r_type,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_header_src,
    output[2:0] io_out_bits_header_dst,
    output[1:0] io_out_bits_payload_addr_beat,
    output[25:0] io_out_bits_payload_addr_block,
    output[5:0] io_out_bits_payload_client_xact_id,
    output io_out_bits_payload_voluntary,
    output[2:0] io_out_bits_payload_r_type,
    output[127:0] io_out_bits_payload_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T202;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T203;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  locked;
  wire T204;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] R41;
  wire[1:0] T205;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[127:0] T45;
  wire[127:0] T46;
  wire[127:0] T47;
  wire T48;
  wire[2:0] T49;
  wire[127:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[5:0] T70;
  wire[5:0] T71;
  wire[5:0] T72;
  wire T73;
  wire[5:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire[25:0] T78;
  wire[25:0] T79;
  wire[25:0] T80;
  wire T81;
  wire[25:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire T97;
  wire[2:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire[2:0] T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire T105;
  wire[2:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R41 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T202 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T203 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T35 & T30;
  assign T30 = T32 | T31;
  assign T31 = 3'h2 == io_out_bits_payload_r_type;
  assign T32 = T34 | T33;
  assign T33 = 3'h1 == io_out_bits_payload_r_type;
  assign T34 = 3'h0 == io_out_bits_payload_r_type;
  assign T35 = io_out_valid & io_out_ready;
  assign T204 = reset ? 1'h0 : T36;
  assign T36 = T43 ? 1'h0 : T37;
  assign T37 = T29 ? T38 : locked;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T40 == 2'h0;
  assign T40 = R41 + 2'h1;
  assign T205 = reset ? 2'h0 : T42;
  assign T42 = T29 ? T40 : R41;
  assign T43 = T35 & T44;
  assign T44 = T30 ^ 1'h1;
  assign io_out_bits_payload_data = T45;
  assign T45 = T53 ? io_in_4_bits_payload_data : T46;
  assign T46 = T52 ? T50 : T47;
  assign T47 = T48 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T48 = T49[1'h0];
  assign T49 = chosen;
  assign T50 = T51 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T51 = T49[1'h0];
  assign T52 = T49[1'h1];
  assign T53 = T49[2'h2];
  assign io_out_bits_payload_r_type = T54;
  assign T54 = T61 ? io_in_4_bits_payload_r_type : T55;
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T57 = T49[1'h0];
  assign T58 = T59 ? io_in_3_bits_payload_r_type : io_in_2_bits_payload_r_type;
  assign T59 = T49[1'h0];
  assign T60 = T49[1'h1];
  assign T61 = T49[2'h2];
  assign io_out_bits_payload_voluntary = T62;
  assign T62 = T69 ? io_in_4_bits_payload_voluntary : T63;
  assign T63 = T68 ? T66 : T64;
  assign T64 = T65 ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign T65 = T49[1'h0];
  assign T66 = T67 ? io_in_3_bits_payload_voluntary : io_in_2_bits_payload_voluntary;
  assign T67 = T49[1'h0];
  assign T68 = T49[1'h1];
  assign T69 = T49[2'h2];
  assign io_out_bits_payload_client_xact_id = T70;
  assign T70 = T77 ? io_in_4_bits_payload_client_xact_id : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T73 = T49[1'h0];
  assign T74 = T75 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T75 = T49[1'h0];
  assign T76 = T49[1'h1];
  assign T77 = T49[2'h2];
  assign io_out_bits_payload_addr_block = T78;
  assign T78 = T85 ? io_in_4_bits_payload_addr_block : T79;
  assign T79 = T84 ? T82 : T80;
  assign T80 = T81 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T81 = T49[1'h0];
  assign T82 = T83 ? io_in_3_bits_payload_addr_block : io_in_2_bits_payload_addr_block;
  assign T83 = T49[1'h0];
  assign T84 = T49[1'h1];
  assign T85 = T49[2'h2];
  assign io_out_bits_payload_addr_beat = T86;
  assign T86 = T93 ? io_in_4_bits_payload_addr_beat : T87;
  assign T87 = T92 ? T90 : T88;
  assign T88 = T89 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T89 = T49[1'h0];
  assign T90 = T91 ? io_in_3_bits_payload_addr_beat : io_in_2_bits_payload_addr_beat;
  assign T91 = T49[1'h0];
  assign T92 = T49[1'h1];
  assign T93 = T49[2'h2];
  assign io_out_bits_header_dst = T94;
  assign T94 = T101 ? io_in_4_bits_header_dst : T95;
  assign T95 = T100 ? T98 : T96;
  assign T96 = T97 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T97 = T49[1'h0];
  assign T98 = T99 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T99 = T49[1'h0];
  assign T100 = T49[1'h1];
  assign T101 = T49[2'h2];
  assign io_out_bits_header_src = T102;
  assign T102 = T109 ? io_in_4_bits_header_src : T103;
  assign T103 = T108 ? T106 : T104;
  assign T104 = T105 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T105 = T49[1'h0];
  assign T106 = T107 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T107 = T49[1'h0];
  assign T108 = T49[1'h1];
  assign T109 = T49[2'h2];
  assign io_out_valid = T110;
  assign T110 = T117 ? io_in_4_valid : T111;
  assign T111 = T116 ? T114 : T112;
  assign T112 = T113 ? io_in_1_valid : io_in_0_valid;
  assign T113 = T49[1'h0];
  assign T114 = T115 ? io_in_3_valid : io_in_2_valid;
  assign T115 = T49[1'h0];
  assign T116 = T49[1'h1];
  assign T117 = T49[2'h2];
  assign io_in_0_ready = T118;
  assign T118 = T119 & io_out_ready;
  assign T119 = locked ? T137 : T120;
  assign T120 = T136 | T121;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T125 | T123;
  assign T123 = io_in_4_valid & T124;
  assign T124 = last_grant < 3'h4;
  assign T125 = T128 | T126;
  assign T126 = io_in_3_valid & T127;
  assign T127 = last_grant < 3'h3;
  assign T128 = T131 | T129;
  assign T129 = io_in_2_valid & T130;
  assign T130 = last_grant < 3'h2;
  assign T131 = T134 | T132;
  assign T132 = io_in_1_valid & T133;
  assign T133 = last_grant < 3'h1;
  assign T134 = io_in_0_valid & T135;
  assign T135 = last_grant < 3'h0;
  assign T136 = last_grant < 3'h0;
  assign T137 = lockIdx == 3'h0;
  assign io_in_1_ready = T138;
  assign T138 = T139 & io_out_ready;
  assign T139 = locked ? T150 : T140;
  assign T140 = T147 | T141;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T143 | io_in_0_valid;
  assign T143 = T144 | T123;
  assign T144 = T145 | T126;
  assign T145 = T146 | T129;
  assign T146 = T134 | T132;
  assign T147 = T149 & T148;
  assign T148 = last_grant < 3'h1;
  assign T149 = T134 ^ 1'h1;
  assign T150 = lockIdx == 3'h1;
  assign io_in_2_ready = T151;
  assign T151 = T152 & io_out_ready;
  assign T152 = locked ? T165 : T153;
  assign T153 = T161 | T154;
  assign T154 = T155 ^ 1'h1;
  assign T155 = T156 | io_in_1_valid;
  assign T156 = T157 | io_in_0_valid;
  assign T157 = T158 | T123;
  assign T158 = T159 | T126;
  assign T159 = T160 | T129;
  assign T160 = T134 | T132;
  assign T161 = T163 & T162;
  assign T162 = last_grant < 3'h2;
  assign T163 = T164 ^ 1'h1;
  assign T164 = T134 | T132;
  assign T165 = lockIdx == 3'h2;
  assign io_in_3_ready = T166;
  assign T166 = T167 & io_out_ready;
  assign T167 = locked ? T182 : T168;
  assign T168 = T177 | T169;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T171 | io_in_2_valid;
  assign T171 = T172 | io_in_1_valid;
  assign T172 = T173 | io_in_0_valid;
  assign T173 = T174 | T123;
  assign T174 = T175 | T126;
  assign T175 = T176 | T129;
  assign T176 = T134 | T132;
  assign T177 = T179 & T178;
  assign T178 = last_grant < 3'h3;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T181 | T129;
  assign T181 = T134 | T132;
  assign T182 = lockIdx == 3'h3;
  assign io_in_4_ready = T183;
  assign T183 = T184 & io_out_ready;
  assign T184 = locked ? T201 : T185;
  assign T185 = T195 | T186;
  assign T186 = T187 ^ 1'h1;
  assign T187 = T188 | io_in_3_valid;
  assign T188 = T189 | io_in_2_valid;
  assign T189 = T190 | io_in_1_valid;
  assign T190 = T191 | io_in_0_valid;
  assign T191 = T192 | T123;
  assign T192 = T193 | T126;
  assign T193 = T194 | T129;
  assign T194 = T134 | T132;
  assign T195 = T197 & T196;
  assign T196 = last_grant < 3'h4;
  assign T197 = T198 ^ 1'h1;
  assign T198 = T199 | T126;
  assign T199 = T200 | T129;
  assign T200 = T134 | T132;
  assign T201 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T43) begin
      locked <= 1'h0;
    end else if(T29) begin
      locked <= T38;
    end
    if(reset) begin
      R41 <= 2'h0;
    end else if(T29) begin
      R41 <= T40;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input  io_in_4_bits_payload_voluntary,
    input [2:0] io_in_4_bits_payload_r_type,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input  io_in_3_bits_payload_voluntary,
    input [2:0] io_in_3_bits_payload_r_type,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input  io_in_2_bits_payload_voluntary,
    input [2:0] io_in_2_bits_payload_r_type,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input  io_in_1_bits_payload_voluntary,
    input [2:0] io_in_1_bits_payload_r_type,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input  io_in_0_bits_payload_voluntary,
    input [2:0] io_in_0_bits_payload_r_type,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_4_ready,
    output io_out_4_valid,
    output[2:0] io_out_4_bits_header_src,
    output[2:0] io_out_4_bits_header_dst,
    output[1:0] io_out_4_bits_payload_addr_beat,
    output[25:0] io_out_4_bits_payload_addr_block,
    output[5:0] io_out_4_bits_payload_client_xact_id,
    output io_out_4_bits_payload_voluntary,
    output[2:0] io_out_4_bits_payload_r_type,
    output[127:0] io_out_4_bits_payload_data,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[2:0] io_out_3_bits_header_src,
    output[2:0] io_out_3_bits_header_dst,
    output[1:0] io_out_3_bits_payload_addr_beat,
    output[25:0] io_out_3_bits_payload_addr_block,
    output[5:0] io_out_3_bits_payload_client_xact_id,
    output io_out_3_bits_payload_voluntary,
    output[2:0] io_out_3_bits_payload_r_type,
    output[127:0] io_out_3_bits_payload_data,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[2:0] io_out_2_bits_header_src,
    output[2:0] io_out_2_bits_header_dst,
    output[1:0] io_out_2_bits_payload_addr_beat,
    output[25:0] io_out_2_bits_payload_addr_block,
    output[5:0] io_out_2_bits_payload_client_xact_id,
    output io_out_2_bits_payload_voluntary,
    output[2:0] io_out_2_bits_payload_r_type,
    output[127:0] io_out_2_bits_payload_data,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[2:0] io_out_1_bits_header_src,
    output[2:0] io_out_1_bits_header_dst,
    output[1:0] io_out_1_bits_payload_addr_beat,
    output[25:0] io_out_1_bits_payload_addr_block,
    output[5:0] io_out_1_bits_payload_client_xact_id,
    output io_out_1_bits_payload_voluntary,
    output[2:0] io_out_1_bits_payload_r_type,
    output[127:0] io_out_1_bits_payload_data,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[2:0] io_out_0_bits_header_src,
    output[2:0] io_out_0_bits_header_dst,
    output[1:0] io_out_0_bits_payload_addr_beat,
    output[25:0] io_out_0_bits_payload_addr_block,
    output[5:0] io_out_0_bits_payload_client_xact_id,
    output io_out_0_bits_payload_voluntary,
    output[2:0] io_out_0_bits_payload_r_type,
    output[127:0] io_out_0_bits_payload_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[2:0] LockingRRArbiter_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_1_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire LockingRRArbiter_2_io_in_4_ready;
  wire LockingRRArbiter_2_io_in_3_ready;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_2_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire LockingRRArbiter_3_io_in_4_ready;
  wire LockingRRArbiter_3_io_in_3_ready;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_3_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire LockingRRArbiter_4_io_in_4_ready;
  wire LockingRRArbiter_4_io_in_3_ready;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr_block;
  wire[5:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_4_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_4_io_out_bits_payload_data;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 3'h4;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 3'h4;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 3'h4;
  assign T6 = io_in_3_valid & T7;
  assign T7 = io_in_3_bits_header_dst == 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = io_in_4_bits_header_dst == 3'h4;
  assign T10 = io_in_0_valid & T11;
  assign T11 = io_in_0_bits_header_dst == 3'h3;
  assign T12 = io_in_1_valid & T13;
  assign T13 = io_in_1_bits_header_dst == 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = io_in_2_bits_header_dst == 3'h3;
  assign T16 = io_in_3_valid & T17;
  assign T17 = io_in_3_bits_header_dst == 3'h3;
  assign T18 = io_in_4_valid & T19;
  assign T19 = io_in_4_bits_header_dst == 3'h3;
  assign T20 = io_in_0_valid & T21;
  assign T21 = io_in_0_bits_header_dst == 3'h2;
  assign T22 = io_in_1_valid & T23;
  assign T23 = io_in_1_bits_header_dst == 3'h2;
  assign T24 = io_in_2_valid & T25;
  assign T25 = io_in_2_bits_header_dst == 3'h2;
  assign T26 = io_in_3_valid & T27;
  assign T27 = io_in_3_bits_header_dst == 3'h2;
  assign T28 = io_in_4_valid & T29;
  assign T29 = io_in_4_bits_header_dst == 3'h2;
  assign T30 = io_in_0_valid & T31;
  assign T31 = io_in_0_bits_header_dst == 3'h1;
  assign T32 = io_in_1_valid & T33;
  assign T33 = io_in_1_bits_header_dst == 3'h1;
  assign T34 = io_in_2_valid & T35;
  assign T35 = io_in_2_bits_header_dst == 3'h1;
  assign T36 = io_in_3_valid & T37;
  assign T37 = io_in_3_bits_header_dst == 3'h1;
  assign T38 = io_in_4_valid & T39;
  assign T39 = io_in_4_bits_header_dst == 3'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = io_in_0_bits_header_dst == 3'h0;
  assign T42 = io_in_1_valid & T43;
  assign T43 = io_in_1_bits_header_dst == 3'h0;
  assign T44 = io_in_2_valid & T45;
  assign T45 = io_in_2_bits_header_dst == 3'h0;
  assign T46 = io_in_3_valid & T47;
  assign T47 = io_in_3_bits_header_dst == 3'h0;
  assign T48 = io_in_4_valid & T49;
  assign T49 = io_in_4_bits_header_dst == 3'h0;
  assign io_out_0_bits_payload_data = LockingRRArbiter_io_out_bits_payload_data;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_voluntary = LockingRRArbiter_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_block = LockingRRArbiter_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_addr_beat = LockingRRArbiter_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_header_dst = LockingRRArbiter_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_io_out_valid;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_1_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_voluntary = LockingRRArbiter_1_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_block = LockingRRArbiter_1_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_addr_beat = LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_2_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_voluntary = LockingRRArbiter_2_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_block = LockingRRArbiter_2_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_addr_beat = LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_out_3_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_3_bits_payload_r_type = LockingRRArbiter_3_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_voluntary = LockingRRArbiter_3_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_block = LockingRRArbiter_3_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_addr_beat = LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_3_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_3_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_4_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_4_bits_payload_r_type = LockingRRArbiter_4_io_out_bits_payload_r_type;
  assign io_out_4_bits_payload_voluntary = LockingRRArbiter_4_io_out_bits_payload_voluntary;
  assign io_out_4_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_addr_block = LockingRRArbiter_4_io_out_bits_payload_addr_block;
  assign io_out_4_bits_payload_addr_beat = LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_4_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_4_valid = LockingRRArbiter_4_io_out_valid;
  assign io_in_0_ready = T50;
  assign T50 = T54 | T51;
  assign T51 = T52;
  assign T52 = LockingRRArbiter_4_io_in_0_ready & T53;
  assign T53 = io_in_0_bits_header_dst == 3'h4;
  assign T54 = T58 | T55;
  assign T55 = T56;
  assign T56 = LockingRRArbiter_3_io_in_0_ready & T57;
  assign T57 = io_in_0_bits_header_dst == 3'h3;
  assign T58 = T62 | T59;
  assign T59 = T60;
  assign T60 = LockingRRArbiter_2_io_in_0_ready & T61;
  assign T61 = io_in_0_bits_header_dst == 3'h2;
  assign T62 = T66 | T63;
  assign T63 = T64;
  assign T64 = LockingRRArbiter_1_io_in_0_ready & T65;
  assign T65 = io_in_0_bits_header_dst == 3'h1;
  assign T66 = T67;
  assign T67 = LockingRRArbiter_io_in_0_ready & T68;
  assign T68 = io_in_0_bits_header_dst == 3'h0;
  assign io_in_1_ready = T69;
  assign T69 = T73 | T70;
  assign T70 = T71;
  assign T71 = LockingRRArbiter_4_io_in_1_ready & T72;
  assign T72 = io_in_1_bits_header_dst == 3'h4;
  assign T73 = T77 | T74;
  assign T74 = T75;
  assign T75 = LockingRRArbiter_3_io_in_1_ready & T76;
  assign T76 = io_in_1_bits_header_dst == 3'h3;
  assign T77 = T81 | T78;
  assign T78 = T79;
  assign T79 = LockingRRArbiter_2_io_in_1_ready & T80;
  assign T80 = io_in_1_bits_header_dst == 3'h2;
  assign T81 = T85 | T82;
  assign T82 = T83;
  assign T83 = LockingRRArbiter_1_io_in_1_ready & T84;
  assign T84 = io_in_1_bits_header_dst == 3'h1;
  assign T85 = T86;
  assign T86 = LockingRRArbiter_io_in_1_ready & T87;
  assign T87 = io_in_1_bits_header_dst == 3'h0;
  assign io_in_2_ready = T88;
  assign T88 = T92 | T89;
  assign T89 = T90;
  assign T90 = LockingRRArbiter_4_io_in_2_ready & T91;
  assign T91 = io_in_2_bits_header_dst == 3'h4;
  assign T92 = T96 | T93;
  assign T93 = T94;
  assign T94 = LockingRRArbiter_3_io_in_2_ready & T95;
  assign T95 = io_in_2_bits_header_dst == 3'h3;
  assign T96 = T100 | T97;
  assign T97 = T98;
  assign T98 = LockingRRArbiter_2_io_in_2_ready & T99;
  assign T99 = io_in_2_bits_header_dst == 3'h2;
  assign T100 = T104 | T101;
  assign T101 = T102;
  assign T102 = LockingRRArbiter_1_io_in_2_ready & T103;
  assign T103 = io_in_2_bits_header_dst == 3'h1;
  assign T104 = T105;
  assign T105 = LockingRRArbiter_io_in_2_ready & T106;
  assign T106 = io_in_2_bits_header_dst == 3'h0;
  assign io_in_3_ready = T107;
  assign T107 = T111 | T108;
  assign T108 = T109;
  assign T109 = LockingRRArbiter_4_io_in_3_ready & T110;
  assign T110 = io_in_3_bits_header_dst == 3'h4;
  assign T111 = T115 | T112;
  assign T112 = T113;
  assign T113 = LockingRRArbiter_3_io_in_3_ready & T114;
  assign T114 = io_in_3_bits_header_dst == 3'h3;
  assign T115 = T119 | T116;
  assign T116 = T117;
  assign T117 = LockingRRArbiter_2_io_in_3_ready & T118;
  assign T118 = io_in_3_bits_header_dst == 3'h2;
  assign T119 = T123 | T120;
  assign T120 = T121;
  assign T121 = LockingRRArbiter_1_io_in_3_ready & T122;
  assign T122 = io_in_3_bits_header_dst == 3'h1;
  assign T123 = T124;
  assign T124 = LockingRRArbiter_io_in_3_ready & T125;
  assign T125 = io_in_3_bits_header_dst == 3'h0;
  assign io_in_4_ready = T126;
  assign T126 = T130 | T127;
  assign T127 = T128;
  assign T128 = LockingRRArbiter_4_io_in_4_ready & T129;
  assign T129 = io_in_4_bits_header_dst == 3'h4;
  assign T130 = T134 | T131;
  assign T131 = T132;
  assign T132 = LockingRRArbiter_3_io_in_4_ready & T133;
  assign T133 = io_in_4_bits_header_dst == 3'h3;
  assign T134 = T138 | T135;
  assign T135 = T136;
  assign T136 = LockingRRArbiter_2_io_in_4_ready & T137;
  assign T137 = io_in_4_bits_header_dst == 3'h2;
  assign T138 = T142 | T139;
  assign T139 = T140;
  assign T140 = LockingRRArbiter_1_io_in_4_ready & T141;
  assign T141 = io_in_4_bits_header_dst == 3'h1;
  assign T142 = T143;
  assign T143 = LockingRRArbiter_io_in_4_ready & T144;
  assign T144 = io_in_4_bits_header_dst == 3'h0;
  LockingRRArbiter_6 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( T48 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_voluntary( io_in_4_bits_payload_voluntary ),
       .io_in_4_bits_payload_r_type( io_in_4_bits_payload_r_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( T46 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_voluntary( io_in_3_bits_payload_voluntary ),
       .io_in_3_bits_payload_r_type( io_in_3_bits_payload_r_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( T44 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( io_in_2_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( T42 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( io_in_1_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( io_in_0_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_6 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( T38 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_voluntary( io_in_4_bits_payload_voluntary ),
       .io_in_4_bits_payload_r_type( io_in_4_bits_payload_r_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( T36 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_voluntary( io_in_3_bits_payload_voluntary ),
       .io_in_3_bits_payload_r_type( io_in_3_bits_payload_r_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T34 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( io_in_2_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T32 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( io_in_1_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T30 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( io_in_0_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_6 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( T28 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_voluntary( io_in_4_bits_payload_voluntary ),
       .io_in_4_bits_payload_r_type( io_in_4_bits_payload_r_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( T26 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_voluntary( io_in_3_bits_payload_voluntary ),
       .io_in_3_bits_payload_r_type( io_in_3_bits_payload_r_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T24 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( io_in_2_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T22 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( io_in_1_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( io_in_0_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_2_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_2_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_2_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_2_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_6 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( T18 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_voluntary( io_in_4_bits_payload_voluntary ),
       .io_in_4_bits_payload_r_type( io_in_4_bits_payload_r_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( T16 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_voluntary( io_in_3_bits_payload_voluntary ),
       .io_in_3_bits_payload_r_type( io_in_3_bits_payload_r_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T14 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( io_in_2_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T12 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( io_in_1_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T10 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( io_in_0_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_3_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_3_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_3_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_3_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_3_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_6 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_4_io_in_4_ready ),
       .io_in_4_valid( T8 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_voluntary( io_in_4_bits_payload_voluntary ),
       .io_in_4_bits_payload_r_type( io_in_4_bits_payload_r_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_4_io_in_3_ready ),
       .io_in_3_valid( T6 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_voluntary( io_in_3_bits_payload_voluntary ),
       .io_in_3_bits_payload_r_type( io_in_3_bits_payload_r_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( io_in_2_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( io_in_1_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( io_in_0_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_4_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_4_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_4_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_4_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_4_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_7(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_header_src,
    output[2:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire T7;
  wire T8;
  reg [2:0] last_grant;
  wire[2:0] T132;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire[2:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire[25:0] T26;
  wire[25:0] T27;
  wire[25:0] T28;
  wire T29;
  wire[25:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire[2:0] T44;
  wire T45;
  wire[2:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T15 ? 3'h1 : T0;
  assign T0 = T13 ? 3'h2 : T1;
  assign T1 = T11 ? 3'h3 : T2;
  assign T2 = T7 ? 3'h4 : T3;
  assign T3 = io_in_0_valid ? 3'h0 : T4;
  assign T4 = io_in_1_valid ? 3'h1 : T5;
  assign T5 = io_in_2_valid ? 3'h2 : T6;
  assign T6 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T7 = io_in_4_valid & T8;
  assign T8 = last_grant < 3'h4;
  assign T132 = reset ? 3'h0 : T9;
  assign T9 = T10 ? chosen : last_grant;
  assign T10 = io_out_ready & io_out_valid;
  assign T11 = io_in_3_valid & T12;
  assign T12 = last_grant < 3'h3;
  assign T13 = io_in_2_valid & T14;
  assign T14 = last_grant < 3'h2;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 3'h1;
  assign io_out_bits_payload_p_type = T17;
  assign T17 = T25 ? io_in_4_bits_payload_p_type : T18;
  assign T18 = T24 ? T22 : T19;
  assign T19 = T20 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T20 = T21[1'h0];
  assign T21 = chosen;
  assign T22 = T23 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T23 = T21[1'h0];
  assign T24 = T21[1'h1];
  assign T25 = T21[2'h2];
  assign io_out_bits_payload_addr_block = T26;
  assign T26 = T33 ? io_in_4_bits_payload_addr_block : T27;
  assign T27 = T32 ? T30 : T28;
  assign T28 = T29 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T29 = T21[1'h0];
  assign T30 = T31 ? io_in_3_bits_payload_addr_block : io_in_2_bits_payload_addr_block;
  assign T31 = T21[1'h0];
  assign T32 = T21[1'h1];
  assign T33 = T21[2'h2];
  assign io_out_bits_header_dst = T34;
  assign T34 = T41 ? io_in_4_bits_header_dst : T35;
  assign T35 = T40 ? T38 : T36;
  assign T36 = T37 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T37 = T21[1'h0];
  assign T38 = T39 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T39 = T21[1'h0];
  assign T40 = T21[1'h1];
  assign T41 = T21[2'h2];
  assign io_out_bits_header_src = T42;
  assign T42 = T49 ? io_in_4_bits_header_src : T43;
  assign T43 = T48 ? T46 : T44;
  assign T44 = T45 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T45 = T21[1'h0];
  assign T46 = T47 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T47 = T21[1'h0];
  assign T48 = T21[1'h1];
  assign T49 = T21[2'h2];
  assign io_out_valid = T50;
  assign T50 = T57 ? io_in_4_valid : T51;
  assign T51 = T56 ? T54 : T52;
  assign T52 = T53 ? io_in_1_valid : io_in_0_valid;
  assign T53 = T21[1'h0];
  assign T54 = T55 ? io_in_3_valid : io_in_2_valid;
  assign T55 = T21[1'h0];
  assign T56 = T21[1'h1];
  assign T57 = T21[2'h2];
  assign io_in_0_ready = T58;
  assign T58 = T59 & io_out_ready;
  assign T59 = T75 | T60;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T64 | T62;
  assign T62 = io_in_4_valid & T63;
  assign T63 = last_grant < 3'h4;
  assign T64 = T67 | T65;
  assign T65 = io_in_3_valid & T66;
  assign T66 = last_grant < 3'h3;
  assign T67 = T70 | T68;
  assign T68 = io_in_2_valid & T69;
  assign T69 = last_grant < 3'h2;
  assign T70 = T73 | T71;
  assign T71 = io_in_1_valid & T72;
  assign T72 = last_grant < 3'h1;
  assign T73 = io_in_0_valid & T74;
  assign T74 = last_grant < 3'h0;
  assign T75 = last_grant < 3'h0;
  assign io_in_1_ready = T76;
  assign T76 = T77 & io_out_ready;
  assign T77 = T84 | T78;
  assign T78 = T79 ^ 1'h1;
  assign T79 = T80 | io_in_0_valid;
  assign T80 = T81 | T62;
  assign T81 = T82 | T65;
  assign T82 = T83 | T68;
  assign T83 = T73 | T71;
  assign T84 = T86 & T85;
  assign T85 = last_grant < 3'h1;
  assign T86 = T73 ^ 1'h1;
  assign io_in_2_ready = T87;
  assign T87 = T88 & io_out_ready;
  assign T88 = T96 | T89;
  assign T89 = T90 ^ 1'h1;
  assign T90 = T91 | io_in_1_valid;
  assign T91 = T92 | io_in_0_valid;
  assign T92 = T93 | T62;
  assign T93 = T94 | T65;
  assign T94 = T95 | T68;
  assign T95 = T73 | T71;
  assign T96 = T98 & T97;
  assign T97 = last_grant < 3'h2;
  assign T98 = T99 ^ 1'h1;
  assign T99 = T73 | T71;
  assign io_in_3_ready = T100;
  assign T100 = T101 & io_out_ready;
  assign T101 = T110 | T102;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T104 | io_in_2_valid;
  assign T104 = T105 | io_in_1_valid;
  assign T105 = T106 | io_in_0_valid;
  assign T106 = T107 | T62;
  assign T107 = T108 | T65;
  assign T108 = T109 | T68;
  assign T109 = T73 | T71;
  assign T110 = T112 & T111;
  assign T111 = last_grant < 3'h3;
  assign T112 = T113 ^ 1'h1;
  assign T113 = T114 | T68;
  assign T114 = T73 | T71;
  assign io_in_4_ready = T115;
  assign T115 = T116 & io_out_ready;
  assign T116 = T126 | T117;
  assign T117 = T118 ^ 1'h1;
  assign T118 = T119 | io_in_3_valid;
  assign T119 = T120 | io_in_2_valid;
  assign T120 = T121 | io_in_1_valid;
  assign T121 = T122 | io_in_0_valid;
  assign T122 = T123 | T62;
  assign T123 = T124 | T65;
  assign T124 = T125 | T68;
  assign T125 = T73 | T71;
  assign T126 = T128 & T127;
  assign T127 = last_grant < 3'h4;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | T65;
  assign T130 = T131 | T68;
  assign T131 = T73 | T71;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T10) begin
      last_grant <= chosen;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr_block,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr_block,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_4_ready,
    output io_out_4_valid,
    output[2:0] io_out_4_bits_header_src,
    output[2:0] io_out_4_bits_header_dst,
    output[25:0] io_out_4_bits_payload_addr_block,
    output[1:0] io_out_4_bits_payload_p_type,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[2:0] io_out_3_bits_header_src,
    output[2:0] io_out_3_bits_header_dst,
    output[25:0] io_out_3_bits_payload_addr_block,
    output[1:0] io_out_3_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[2:0] io_out_2_bits_header_src,
    output[2:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr_block,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[2:0] io_out_1_bits_header_src,
    output[2:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr_block,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[2:0] io_out_0_bits_header_src,
    output[2:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr_block,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[2:0] LockingRRArbiter_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_p_type;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_p_type;
  wire LockingRRArbiter_2_io_in_4_ready;
  wire LockingRRArbiter_2_io_in_3_ready;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_p_type;
  wire LockingRRArbiter_3_io_in_4_ready;
  wire LockingRRArbiter_3_io_in_3_ready;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_p_type;
  wire LockingRRArbiter_4_io_in_4_ready;
  wire LockingRRArbiter_4_io_in_3_ready;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_p_type;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 3'h4;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 3'h4;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 3'h4;
  assign T6 = io_in_3_valid & T7;
  assign T7 = io_in_3_bits_header_dst == 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = io_in_4_bits_header_dst == 3'h4;
  assign T10 = io_in_0_valid & T11;
  assign T11 = io_in_0_bits_header_dst == 3'h3;
  assign T12 = io_in_1_valid & T13;
  assign T13 = io_in_1_bits_header_dst == 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = io_in_2_bits_header_dst == 3'h3;
  assign T16 = io_in_3_valid & T17;
  assign T17 = io_in_3_bits_header_dst == 3'h3;
  assign T18 = io_in_4_valid & T19;
  assign T19 = io_in_4_bits_header_dst == 3'h3;
  assign T20 = io_in_0_valid & T21;
  assign T21 = io_in_0_bits_header_dst == 3'h2;
  assign T22 = io_in_1_valid & T23;
  assign T23 = io_in_1_bits_header_dst == 3'h2;
  assign T24 = io_in_2_valid & T25;
  assign T25 = io_in_2_bits_header_dst == 3'h2;
  assign T26 = io_in_3_valid & T27;
  assign T27 = io_in_3_bits_header_dst == 3'h2;
  assign T28 = io_in_4_valid & T29;
  assign T29 = io_in_4_bits_header_dst == 3'h2;
  assign T30 = io_in_0_valid & T31;
  assign T31 = io_in_0_bits_header_dst == 3'h1;
  assign T32 = io_in_1_valid & T33;
  assign T33 = io_in_1_bits_header_dst == 3'h1;
  assign T34 = io_in_2_valid & T35;
  assign T35 = io_in_2_bits_header_dst == 3'h1;
  assign T36 = io_in_3_valid & T37;
  assign T37 = io_in_3_bits_header_dst == 3'h1;
  assign T38 = io_in_4_valid & T39;
  assign T39 = io_in_4_bits_header_dst == 3'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = io_in_0_bits_header_dst == 3'h0;
  assign T42 = io_in_1_valid & T43;
  assign T43 = io_in_1_bits_header_dst == 3'h0;
  assign T44 = io_in_2_valid & T45;
  assign T45 = io_in_2_bits_header_dst == 3'h0;
  assign T46 = io_in_3_valid & T47;
  assign T47 = io_in_3_bits_header_dst == 3'h0;
  assign T48 = io_in_4_valid & T49;
  assign T49 = io_in_4_bits_header_dst == 3'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_addr_block = LockingRRArbiter_io_out_bits_payload_addr_block;
  assign io_out_0_bits_header_dst = LockingRRArbiter_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_1_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_addr_block = LockingRRArbiter_1_io_out_bits_payload_addr_block;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_2_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_addr_block = LockingRRArbiter_2_io_out_bits_payload_addr_block;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_out_3_bits_payload_p_type = LockingRRArbiter_3_io_out_bits_payload_p_type;
  assign io_out_3_bits_payload_addr_block = LockingRRArbiter_3_io_out_bits_payload_addr_block;
  assign io_out_3_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_3_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_3_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_4_bits_payload_p_type = LockingRRArbiter_4_io_out_bits_payload_p_type;
  assign io_out_4_bits_payload_addr_block = LockingRRArbiter_4_io_out_bits_payload_addr_block;
  assign io_out_4_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_4_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_4_valid = LockingRRArbiter_4_io_out_valid;
  assign io_in_0_ready = T50;
  assign T50 = T54 | T51;
  assign T51 = T52;
  assign T52 = LockingRRArbiter_4_io_in_0_ready & T53;
  assign T53 = io_in_0_bits_header_dst == 3'h4;
  assign T54 = T58 | T55;
  assign T55 = T56;
  assign T56 = LockingRRArbiter_3_io_in_0_ready & T57;
  assign T57 = io_in_0_bits_header_dst == 3'h3;
  assign T58 = T62 | T59;
  assign T59 = T60;
  assign T60 = LockingRRArbiter_2_io_in_0_ready & T61;
  assign T61 = io_in_0_bits_header_dst == 3'h2;
  assign T62 = T66 | T63;
  assign T63 = T64;
  assign T64 = LockingRRArbiter_1_io_in_0_ready & T65;
  assign T65 = io_in_0_bits_header_dst == 3'h1;
  assign T66 = T67;
  assign T67 = LockingRRArbiter_io_in_0_ready & T68;
  assign T68 = io_in_0_bits_header_dst == 3'h0;
  assign io_in_1_ready = T69;
  assign T69 = T73 | T70;
  assign T70 = T71;
  assign T71 = LockingRRArbiter_4_io_in_1_ready & T72;
  assign T72 = io_in_1_bits_header_dst == 3'h4;
  assign T73 = T77 | T74;
  assign T74 = T75;
  assign T75 = LockingRRArbiter_3_io_in_1_ready & T76;
  assign T76 = io_in_1_bits_header_dst == 3'h3;
  assign T77 = T81 | T78;
  assign T78 = T79;
  assign T79 = LockingRRArbiter_2_io_in_1_ready & T80;
  assign T80 = io_in_1_bits_header_dst == 3'h2;
  assign T81 = T85 | T82;
  assign T82 = T83;
  assign T83 = LockingRRArbiter_1_io_in_1_ready & T84;
  assign T84 = io_in_1_bits_header_dst == 3'h1;
  assign T85 = T86;
  assign T86 = LockingRRArbiter_io_in_1_ready & T87;
  assign T87 = io_in_1_bits_header_dst == 3'h0;
  assign io_in_2_ready = T88;
  assign T88 = T92 | T89;
  assign T89 = T90;
  assign T90 = LockingRRArbiter_4_io_in_2_ready & T91;
  assign T91 = io_in_2_bits_header_dst == 3'h4;
  assign T92 = T96 | T93;
  assign T93 = T94;
  assign T94 = LockingRRArbiter_3_io_in_2_ready & T95;
  assign T95 = io_in_2_bits_header_dst == 3'h3;
  assign T96 = T100 | T97;
  assign T97 = T98;
  assign T98 = LockingRRArbiter_2_io_in_2_ready & T99;
  assign T99 = io_in_2_bits_header_dst == 3'h2;
  assign T100 = T104 | T101;
  assign T101 = T102;
  assign T102 = LockingRRArbiter_1_io_in_2_ready & T103;
  assign T103 = io_in_2_bits_header_dst == 3'h1;
  assign T104 = T105;
  assign T105 = LockingRRArbiter_io_in_2_ready & T106;
  assign T106 = io_in_2_bits_header_dst == 3'h0;
  assign io_in_3_ready = T107;
  assign T107 = T111 | T108;
  assign T108 = T109;
  assign T109 = LockingRRArbiter_4_io_in_3_ready & T110;
  assign T110 = io_in_3_bits_header_dst == 3'h4;
  assign T111 = T115 | T112;
  assign T112 = T113;
  assign T113 = LockingRRArbiter_3_io_in_3_ready & T114;
  assign T114 = io_in_3_bits_header_dst == 3'h3;
  assign T115 = T119 | T116;
  assign T116 = T117;
  assign T117 = LockingRRArbiter_2_io_in_3_ready & T118;
  assign T118 = io_in_3_bits_header_dst == 3'h2;
  assign T119 = T123 | T120;
  assign T120 = T121;
  assign T121 = LockingRRArbiter_1_io_in_3_ready & T122;
  assign T122 = io_in_3_bits_header_dst == 3'h1;
  assign T123 = T124;
  assign T124 = LockingRRArbiter_io_in_3_ready & T125;
  assign T125 = io_in_3_bits_header_dst == 3'h0;
  assign io_in_4_ready = T126;
  assign T126 = T130 | T127;
  assign T127 = T128;
  assign T128 = LockingRRArbiter_4_io_in_4_ready & T129;
  assign T129 = io_in_4_bits_header_dst == 3'h4;
  assign T130 = T134 | T131;
  assign T131 = T132;
  assign T132 = LockingRRArbiter_3_io_in_4_ready & T133;
  assign T133 = io_in_4_bits_header_dst == 3'h3;
  assign T134 = T138 | T135;
  assign T135 = T136;
  assign T136 = LockingRRArbiter_2_io_in_4_ready & T137;
  assign T137 = io_in_4_bits_header_dst == 3'h2;
  assign T138 = T142 | T139;
  assign T139 = T140;
  assign T140 = LockingRRArbiter_1_io_in_4_ready & T141;
  assign T141 = io_in_4_bits_header_dst == 3'h1;
  assign T142 = T143;
  assign T143 = LockingRRArbiter_io_in_4_ready & T144;
  assign T144 = io_in_4_bits_header_dst == 3'h0;
  LockingRRArbiter_7 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( T48 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_p_type( io_in_4_bits_payload_p_type ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( T46 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_p_type( io_in_3_bits_payload_p_type ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( T44 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( T42 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_p_type( LockingRRArbiter_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_7 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( T38 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_p_type( io_in_4_bits_payload_p_type ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( T36 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_p_type( io_in_3_bits_payload_p_type ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T34 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T32 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T30 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_p_type( LockingRRArbiter_1_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_7 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( T28 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_p_type( io_in_4_bits_payload_p_type ),
       .io_in_3_ready( LockingRRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( T26 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_p_type( io_in_3_bits_payload_p_type ),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T24 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T22 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_2_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_p_type( LockingRRArbiter_2_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_7 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( T18 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_p_type( io_in_4_bits_payload_p_type ),
       .io_in_3_ready( LockingRRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( T16 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_p_type( io_in_3_bits_payload_p_type ),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T14 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T12 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T10 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_3_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_3_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_p_type( LockingRRArbiter_3_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_7 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_4_io_in_4_ready ),
       .io_in_4_valid( T8 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_block( io_in_4_bits_payload_addr_block ),
       .io_in_4_bits_payload_p_type( io_in_4_bits_payload_p_type ),
       .io_in_3_ready( LockingRRArbiter_4_io_in_3_ready ),
       .io_in_3_valid( T6 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_block( io_in_3_bits_payload_addr_block ),
       .io_in_3_bits_payload_p_type( io_in_3_bits_payload_p_type ),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( io_in_2_bits_payload_addr_block ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( io_in_1_bits_payload_addr_block ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( io_in_0_bits_payload_addr_block ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_4_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_4_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_p_type( LockingRRArbiter_4_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_8(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input [3:0] io_in_4_bits_payload_manager_xact_id,
    input  io_in_4_bits_payload_is_builtin_type,
    input [3:0] io_in_4_bits_payload_g_type,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input [3:0] io_in_3_bits_payload_manager_xact_id,
    input  io_in_3_bits_payload_is_builtin_type,
    input [3:0] io_in_3_bits_payload_g_type,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    input  io_in_2_bits_payload_is_builtin_type,
    input [3:0] io_in_2_bits_payload_g_type,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    input  io_in_1_bits_payload_is_builtin_type,
    input [3:0] io_in_1_bits_payload_g_type,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_is_builtin_type,
    input [3:0] io_in_0_bits_payload_g_type,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_header_src,
    output[2:0] io_out_bits_header_dst,
    output[1:0] io_out_bits_payload_addr_beat,
    output[5:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_out_bits_payload_is_builtin_type,
    output[3:0] io_out_bits_payload_g_type,
    output[127:0] io_out_bits_payload_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T202;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T203;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  locked;
  wire T204;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] R41;
  wire[1:0] T205;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[127:0] T45;
  wire[127:0] T46;
  wire[127:0] T47;
  wire T48;
  wire[2:0] T49;
  wire[127:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[3:0] T56;
  wire T57;
  wire[3:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire T73;
  wire[3:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire[5:0] T78;
  wire[5:0] T79;
  wire[5:0] T80;
  wire T81;
  wire[5:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire T97;
  wire[2:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire[2:0] T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire T105;
  wire[2:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R41 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T202 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T203 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T35 & T30;
  assign T30 = io_out_bits_payload_is_builtin_type ? T34 : T31;
  assign T31 = T33 | T32;
  assign T32 = 4'h1 == io_out_bits_payload_g_type;
  assign T33 = 4'h0 == io_out_bits_payload_g_type;
  assign T34 = 4'h5 == io_out_bits_payload_g_type;
  assign T35 = io_out_valid & io_out_ready;
  assign T204 = reset ? 1'h0 : T36;
  assign T36 = T43 ? 1'h0 : T37;
  assign T37 = T29 ? T38 : locked;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T40 == 2'h0;
  assign T40 = R41 + 2'h1;
  assign T205 = reset ? 2'h0 : T42;
  assign T42 = T29 ? T40 : R41;
  assign T43 = T35 & T44;
  assign T44 = T30 ^ 1'h1;
  assign io_out_bits_payload_data = T45;
  assign T45 = T53 ? io_in_4_bits_payload_data : T46;
  assign T46 = T52 ? T50 : T47;
  assign T47 = T48 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T48 = T49[1'h0];
  assign T49 = chosen;
  assign T50 = T51 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T51 = T49[1'h0];
  assign T52 = T49[1'h1];
  assign T53 = T49[2'h2];
  assign io_out_bits_payload_g_type = T54;
  assign T54 = T61 ? io_in_4_bits_payload_g_type : T55;
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T57 = T49[1'h0];
  assign T58 = T59 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T59 = T49[1'h0];
  assign T60 = T49[1'h1];
  assign T61 = T49[2'h2];
  assign io_out_bits_payload_is_builtin_type = T62;
  assign T62 = T69 ? io_in_4_bits_payload_is_builtin_type : T63;
  assign T63 = T68 ? T66 : T64;
  assign T64 = T65 ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign T65 = T49[1'h0];
  assign T66 = T67 ? io_in_3_bits_payload_is_builtin_type : io_in_2_bits_payload_is_builtin_type;
  assign T67 = T49[1'h0];
  assign T68 = T49[1'h1];
  assign T69 = T49[2'h2];
  assign io_out_bits_payload_manager_xact_id = T70;
  assign T70 = T77 ? io_in_4_bits_payload_manager_xact_id : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T73 = T49[1'h0];
  assign T74 = T75 ? io_in_3_bits_payload_manager_xact_id : io_in_2_bits_payload_manager_xact_id;
  assign T75 = T49[1'h0];
  assign T76 = T49[1'h1];
  assign T77 = T49[2'h2];
  assign io_out_bits_payload_client_xact_id = T78;
  assign T78 = T85 ? io_in_4_bits_payload_client_xact_id : T79;
  assign T79 = T84 ? T82 : T80;
  assign T80 = T81 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T81 = T49[1'h0];
  assign T82 = T83 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T83 = T49[1'h0];
  assign T84 = T49[1'h1];
  assign T85 = T49[2'h2];
  assign io_out_bits_payload_addr_beat = T86;
  assign T86 = T93 ? io_in_4_bits_payload_addr_beat : T87;
  assign T87 = T92 ? T90 : T88;
  assign T88 = T89 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T89 = T49[1'h0];
  assign T90 = T91 ? io_in_3_bits_payload_addr_beat : io_in_2_bits_payload_addr_beat;
  assign T91 = T49[1'h0];
  assign T92 = T49[1'h1];
  assign T93 = T49[2'h2];
  assign io_out_bits_header_dst = T94;
  assign T94 = T101 ? io_in_4_bits_header_dst : T95;
  assign T95 = T100 ? T98 : T96;
  assign T96 = T97 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T97 = T49[1'h0];
  assign T98 = T99 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T99 = T49[1'h0];
  assign T100 = T49[1'h1];
  assign T101 = T49[2'h2];
  assign io_out_bits_header_src = T102;
  assign T102 = T109 ? io_in_4_bits_header_src : T103;
  assign T103 = T108 ? T106 : T104;
  assign T104 = T105 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T105 = T49[1'h0];
  assign T106 = T107 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T107 = T49[1'h0];
  assign T108 = T49[1'h1];
  assign T109 = T49[2'h2];
  assign io_out_valid = T110;
  assign T110 = T117 ? io_in_4_valid : T111;
  assign T111 = T116 ? T114 : T112;
  assign T112 = T113 ? io_in_1_valid : io_in_0_valid;
  assign T113 = T49[1'h0];
  assign T114 = T115 ? io_in_3_valid : io_in_2_valid;
  assign T115 = T49[1'h0];
  assign T116 = T49[1'h1];
  assign T117 = T49[2'h2];
  assign io_in_0_ready = T118;
  assign T118 = T119 & io_out_ready;
  assign T119 = locked ? T137 : T120;
  assign T120 = T136 | T121;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T125 | T123;
  assign T123 = io_in_4_valid & T124;
  assign T124 = last_grant < 3'h4;
  assign T125 = T128 | T126;
  assign T126 = io_in_3_valid & T127;
  assign T127 = last_grant < 3'h3;
  assign T128 = T131 | T129;
  assign T129 = io_in_2_valid & T130;
  assign T130 = last_grant < 3'h2;
  assign T131 = T134 | T132;
  assign T132 = io_in_1_valid & T133;
  assign T133 = last_grant < 3'h1;
  assign T134 = io_in_0_valid & T135;
  assign T135 = last_grant < 3'h0;
  assign T136 = last_grant < 3'h0;
  assign T137 = lockIdx == 3'h0;
  assign io_in_1_ready = T138;
  assign T138 = T139 & io_out_ready;
  assign T139 = locked ? T150 : T140;
  assign T140 = T147 | T141;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T143 | io_in_0_valid;
  assign T143 = T144 | T123;
  assign T144 = T145 | T126;
  assign T145 = T146 | T129;
  assign T146 = T134 | T132;
  assign T147 = T149 & T148;
  assign T148 = last_grant < 3'h1;
  assign T149 = T134 ^ 1'h1;
  assign T150 = lockIdx == 3'h1;
  assign io_in_2_ready = T151;
  assign T151 = T152 & io_out_ready;
  assign T152 = locked ? T165 : T153;
  assign T153 = T161 | T154;
  assign T154 = T155 ^ 1'h1;
  assign T155 = T156 | io_in_1_valid;
  assign T156 = T157 | io_in_0_valid;
  assign T157 = T158 | T123;
  assign T158 = T159 | T126;
  assign T159 = T160 | T129;
  assign T160 = T134 | T132;
  assign T161 = T163 & T162;
  assign T162 = last_grant < 3'h2;
  assign T163 = T164 ^ 1'h1;
  assign T164 = T134 | T132;
  assign T165 = lockIdx == 3'h2;
  assign io_in_3_ready = T166;
  assign T166 = T167 & io_out_ready;
  assign T167 = locked ? T182 : T168;
  assign T168 = T177 | T169;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T171 | io_in_2_valid;
  assign T171 = T172 | io_in_1_valid;
  assign T172 = T173 | io_in_0_valid;
  assign T173 = T174 | T123;
  assign T174 = T175 | T126;
  assign T175 = T176 | T129;
  assign T176 = T134 | T132;
  assign T177 = T179 & T178;
  assign T178 = last_grant < 3'h3;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T181 | T129;
  assign T181 = T134 | T132;
  assign T182 = lockIdx == 3'h3;
  assign io_in_4_ready = T183;
  assign T183 = T184 & io_out_ready;
  assign T184 = locked ? T201 : T185;
  assign T185 = T195 | T186;
  assign T186 = T187 ^ 1'h1;
  assign T187 = T188 | io_in_3_valid;
  assign T188 = T189 | io_in_2_valid;
  assign T189 = T190 | io_in_1_valid;
  assign T190 = T191 | io_in_0_valid;
  assign T191 = T192 | T123;
  assign T192 = T193 | T126;
  assign T193 = T194 | T129;
  assign T194 = T134 | T132;
  assign T195 = T197 & T196;
  assign T196 = last_grant < 3'h4;
  assign T197 = T198 ^ 1'h1;
  assign T198 = T199 | T126;
  assign T199 = T200 | T129;
  assign T200 = T134 | T132;
  assign T201 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T43) begin
      locked <= 1'h0;
    end else if(T29) begin
      locked <= T38;
    end
    if(reset) begin
      R41 <= 2'h0;
    end else if(T29) begin
      R41 <= T40;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [1:0] io_in_4_bits_payload_addr_beat,
    input [5:0] io_in_4_bits_payload_client_xact_id,
    input [3:0] io_in_4_bits_payload_manager_xact_id,
    input  io_in_4_bits_payload_is_builtin_type,
    input [3:0] io_in_4_bits_payload_g_type,
    input [127:0] io_in_4_bits_payload_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [1:0] io_in_3_bits_payload_addr_beat,
    input [5:0] io_in_3_bits_payload_client_xact_id,
    input [3:0] io_in_3_bits_payload_manager_xact_id,
    input  io_in_3_bits_payload_is_builtin_type,
    input [3:0] io_in_3_bits_payload_g_type,
    input [127:0] io_in_3_bits_payload_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [5:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    input  io_in_2_bits_payload_is_builtin_type,
    input [3:0] io_in_2_bits_payload_g_type,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [5:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    input  io_in_1_bits_payload_is_builtin_type,
    input [3:0] io_in_1_bits_payload_g_type,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [5:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_is_builtin_type,
    input [3:0] io_in_0_bits_payload_g_type,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_4_ready,
    output io_out_4_valid,
    output[2:0] io_out_4_bits_header_src,
    output[2:0] io_out_4_bits_header_dst,
    output[1:0] io_out_4_bits_payload_addr_beat,
    output[5:0] io_out_4_bits_payload_client_xact_id,
    output[3:0] io_out_4_bits_payload_manager_xact_id,
    output io_out_4_bits_payload_is_builtin_type,
    output[3:0] io_out_4_bits_payload_g_type,
    output[127:0] io_out_4_bits_payload_data,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[2:0] io_out_3_bits_header_src,
    output[2:0] io_out_3_bits_header_dst,
    output[1:0] io_out_3_bits_payload_addr_beat,
    output[5:0] io_out_3_bits_payload_client_xact_id,
    output[3:0] io_out_3_bits_payload_manager_xact_id,
    output io_out_3_bits_payload_is_builtin_type,
    output[3:0] io_out_3_bits_payload_g_type,
    output[127:0] io_out_3_bits_payload_data,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[2:0] io_out_2_bits_header_src,
    output[2:0] io_out_2_bits_header_dst,
    output[1:0] io_out_2_bits_payload_addr_beat,
    output[5:0] io_out_2_bits_payload_client_xact_id,
    output[3:0] io_out_2_bits_payload_manager_xact_id,
    output io_out_2_bits_payload_is_builtin_type,
    output[3:0] io_out_2_bits_payload_g_type,
    output[127:0] io_out_2_bits_payload_data,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[2:0] io_out_1_bits_header_src,
    output[2:0] io_out_1_bits_header_dst,
    output[1:0] io_out_1_bits_payload_addr_beat,
    output[5:0] io_out_1_bits_payload_client_xact_id,
    output[3:0] io_out_1_bits_payload_manager_xact_id,
    output io_out_1_bits_payload_is_builtin_type,
    output[3:0] io_out_1_bits_payload_g_type,
    output[127:0] io_out_1_bits_payload_data,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[2:0] io_out_0_bits_header_src,
    output[2:0] io_out_0_bits_header_dst,
    output[1:0] io_out_0_bits_payload_addr_beat,
    output[5:0] io_out_0_bits_payload_client_xact_id,
    output[3:0] io_out_0_bits_payload_manager_xact_id,
    output io_out_0_bits_payload_is_builtin_type,
    output[3:0] io_out_0_bits_payload_g_type,
    output[127:0] io_out_0_bits_payload_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[2:0] LockingRRArbiter_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire[5:0] LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  wire[3:0] LockingRRArbiter_io_out_bits_payload_g_type;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_1_io_out_bits_payload_is_builtin_type;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_g_type;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire LockingRRArbiter_2_io_in_4_ready;
  wire LockingRRArbiter_2_io_in_3_ready;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_2_io_out_bits_payload_is_builtin_type;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_g_type;
  wire[127:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire LockingRRArbiter_3_io_in_4_ready;
  wire LockingRRArbiter_3_io_in_3_ready;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  wire[5:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_3_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_3_io_out_bits_payload_is_builtin_type;
  wire[3:0] LockingRRArbiter_3_io_out_bits_payload_g_type;
  wire[127:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire LockingRRArbiter_4_io_in_4_ready;
  wire LockingRRArbiter_4_io_in_3_ready;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  wire[5:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_4_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_4_io_out_bits_payload_is_builtin_type;
  wire[3:0] LockingRRArbiter_4_io_out_bits_payload_g_type;
  wire[127:0] LockingRRArbiter_4_io_out_bits_payload_data;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 3'h4;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 3'h4;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 3'h4;
  assign T6 = io_in_3_valid & T7;
  assign T7 = io_in_3_bits_header_dst == 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = io_in_4_bits_header_dst == 3'h4;
  assign T10 = io_in_0_valid & T11;
  assign T11 = io_in_0_bits_header_dst == 3'h3;
  assign T12 = io_in_1_valid & T13;
  assign T13 = io_in_1_bits_header_dst == 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = io_in_2_bits_header_dst == 3'h3;
  assign T16 = io_in_3_valid & T17;
  assign T17 = io_in_3_bits_header_dst == 3'h3;
  assign T18 = io_in_4_valid & T19;
  assign T19 = io_in_4_bits_header_dst == 3'h3;
  assign T20 = io_in_0_valid & T21;
  assign T21 = io_in_0_bits_header_dst == 3'h2;
  assign T22 = io_in_1_valid & T23;
  assign T23 = io_in_1_bits_header_dst == 3'h2;
  assign T24 = io_in_2_valid & T25;
  assign T25 = io_in_2_bits_header_dst == 3'h2;
  assign T26 = io_in_3_valid & T27;
  assign T27 = io_in_3_bits_header_dst == 3'h2;
  assign T28 = io_in_4_valid & T29;
  assign T29 = io_in_4_bits_header_dst == 3'h2;
  assign T30 = io_in_0_valid & T31;
  assign T31 = io_in_0_bits_header_dst == 3'h1;
  assign T32 = io_in_1_valid & T33;
  assign T33 = io_in_1_bits_header_dst == 3'h1;
  assign T34 = io_in_2_valid & T35;
  assign T35 = io_in_2_bits_header_dst == 3'h1;
  assign T36 = io_in_3_valid & T37;
  assign T37 = io_in_3_bits_header_dst == 3'h1;
  assign T38 = io_in_4_valid & T39;
  assign T39 = io_in_4_bits_header_dst == 3'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = io_in_0_bits_header_dst == 3'h0;
  assign T42 = io_in_1_valid & T43;
  assign T43 = io_in_1_bits_header_dst == 3'h0;
  assign T44 = io_in_2_valid & T45;
  assign T45 = io_in_2_bits_header_dst == 3'h0;
  assign T46 = io_in_3_valid & T47;
  assign T47 = io_in_3_bits_header_dst == 3'h0;
  assign T48 = io_in_4_valid & T49;
  assign T49 = io_in_4_bits_header_dst == 3'h0;
  assign io_out_0_bits_payload_data = LockingRRArbiter_io_out_bits_payload_data;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_is_builtin_type = LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_manager_xact_id = LockingRRArbiter_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = LockingRRArbiter_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_header_dst = LockingRRArbiter_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_io_out_valid;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_1_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_is_builtin_type = LockingRRArbiter_1_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_manager_xact_id = LockingRRArbiter_1_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_2_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_is_builtin_type = LockingRRArbiter_2_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_manager_xact_id = LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = LockingRRArbiter_2_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_out_3_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_3_bits_payload_g_type = LockingRRArbiter_3_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_is_builtin_type = LockingRRArbiter_3_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_manager_xact_id = LockingRRArbiter_3_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = LockingRRArbiter_3_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_3_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_3_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_4_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_4_bits_payload_g_type = LockingRRArbiter_4_io_out_bits_payload_g_type;
  assign io_out_4_bits_payload_is_builtin_type = LockingRRArbiter_4_io_out_bits_payload_is_builtin_type;
  assign io_out_4_bits_payload_manager_xact_id = LockingRRArbiter_4_io_out_bits_payload_manager_xact_id;
  assign io_out_4_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_addr_beat = LockingRRArbiter_4_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_4_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_4_valid = LockingRRArbiter_4_io_out_valid;
  assign io_in_0_ready = T50;
  assign T50 = T54 | T51;
  assign T51 = T52;
  assign T52 = LockingRRArbiter_4_io_in_0_ready & T53;
  assign T53 = io_in_0_bits_header_dst == 3'h4;
  assign T54 = T58 | T55;
  assign T55 = T56;
  assign T56 = LockingRRArbiter_3_io_in_0_ready & T57;
  assign T57 = io_in_0_bits_header_dst == 3'h3;
  assign T58 = T62 | T59;
  assign T59 = T60;
  assign T60 = LockingRRArbiter_2_io_in_0_ready & T61;
  assign T61 = io_in_0_bits_header_dst == 3'h2;
  assign T62 = T66 | T63;
  assign T63 = T64;
  assign T64 = LockingRRArbiter_1_io_in_0_ready & T65;
  assign T65 = io_in_0_bits_header_dst == 3'h1;
  assign T66 = T67;
  assign T67 = LockingRRArbiter_io_in_0_ready & T68;
  assign T68 = io_in_0_bits_header_dst == 3'h0;
  assign io_in_1_ready = T69;
  assign T69 = T73 | T70;
  assign T70 = T71;
  assign T71 = LockingRRArbiter_4_io_in_1_ready & T72;
  assign T72 = io_in_1_bits_header_dst == 3'h4;
  assign T73 = T77 | T74;
  assign T74 = T75;
  assign T75 = LockingRRArbiter_3_io_in_1_ready & T76;
  assign T76 = io_in_1_bits_header_dst == 3'h3;
  assign T77 = T81 | T78;
  assign T78 = T79;
  assign T79 = LockingRRArbiter_2_io_in_1_ready & T80;
  assign T80 = io_in_1_bits_header_dst == 3'h2;
  assign T81 = T85 | T82;
  assign T82 = T83;
  assign T83 = LockingRRArbiter_1_io_in_1_ready & T84;
  assign T84 = io_in_1_bits_header_dst == 3'h1;
  assign T85 = T86;
  assign T86 = LockingRRArbiter_io_in_1_ready & T87;
  assign T87 = io_in_1_bits_header_dst == 3'h0;
  assign io_in_2_ready = T88;
  assign T88 = T92 | T89;
  assign T89 = T90;
  assign T90 = LockingRRArbiter_4_io_in_2_ready & T91;
  assign T91 = io_in_2_bits_header_dst == 3'h4;
  assign T92 = T96 | T93;
  assign T93 = T94;
  assign T94 = LockingRRArbiter_3_io_in_2_ready & T95;
  assign T95 = io_in_2_bits_header_dst == 3'h3;
  assign T96 = T100 | T97;
  assign T97 = T98;
  assign T98 = LockingRRArbiter_2_io_in_2_ready & T99;
  assign T99 = io_in_2_bits_header_dst == 3'h2;
  assign T100 = T104 | T101;
  assign T101 = T102;
  assign T102 = LockingRRArbiter_1_io_in_2_ready & T103;
  assign T103 = io_in_2_bits_header_dst == 3'h1;
  assign T104 = T105;
  assign T105 = LockingRRArbiter_io_in_2_ready & T106;
  assign T106 = io_in_2_bits_header_dst == 3'h0;
  assign io_in_3_ready = T107;
  assign T107 = T111 | T108;
  assign T108 = T109;
  assign T109 = LockingRRArbiter_4_io_in_3_ready & T110;
  assign T110 = io_in_3_bits_header_dst == 3'h4;
  assign T111 = T115 | T112;
  assign T112 = T113;
  assign T113 = LockingRRArbiter_3_io_in_3_ready & T114;
  assign T114 = io_in_3_bits_header_dst == 3'h3;
  assign T115 = T119 | T116;
  assign T116 = T117;
  assign T117 = LockingRRArbiter_2_io_in_3_ready & T118;
  assign T118 = io_in_3_bits_header_dst == 3'h2;
  assign T119 = T123 | T120;
  assign T120 = T121;
  assign T121 = LockingRRArbiter_1_io_in_3_ready & T122;
  assign T122 = io_in_3_bits_header_dst == 3'h1;
  assign T123 = T124;
  assign T124 = LockingRRArbiter_io_in_3_ready & T125;
  assign T125 = io_in_3_bits_header_dst == 3'h0;
  assign io_in_4_ready = T126;
  assign T126 = T130 | T127;
  assign T127 = T128;
  assign T128 = LockingRRArbiter_4_io_in_4_ready & T129;
  assign T129 = io_in_4_bits_header_dst == 3'h4;
  assign T130 = T134 | T131;
  assign T131 = T132;
  assign T132 = LockingRRArbiter_3_io_in_4_ready & T133;
  assign T133 = io_in_4_bits_header_dst == 3'h3;
  assign T134 = T138 | T135;
  assign T135 = T136;
  assign T136 = LockingRRArbiter_2_io_in_4_ready & T137;
  assign T137 = io_in_4_bits_header_dst == 3'h2;
  assign T138 = T142 | T139;
  assign T139 = T140;
  assign T140 = LockingRRArbiter_1_io_in_4_ready & T141;
  assign T141 = io_in_4_bits_header_dst == 3'h1;
  assign T142 = T143;
  assign T143 = LockingRRArbiter_io_in_4_ready & T144;
  assign T144 = io_in_4_bits_header_dst == 3'h0;
  LockingRRArbiter_8 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( T48 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_g_type( io_in_4_bits_payload_g_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( T46 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_g_type( io_in_3_bits_payload_g_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( T44 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( T42 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_g_type( LockingRRArbiter_io_out_bits_payload_g_type ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_8 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( T38 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_g_type( io_in_4_bits_payload_g_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( T36 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_g_type( io_in_3_bits_payload_g_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T34 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T32 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T30 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_1_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_1_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_g_type( LockingRRArbiter_1_io_out_bits_payload_g_type ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_8 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( T28 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_g_type( io_in_4_bits_payload_g_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( T26 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_g_type( io_in_3_bits_payload_g_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T24 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T22 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_2_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_2_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_2_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_g_type( LockingRRArbiter_2_io_out_bits_payload_g_type ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_8 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( T18 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_g_type( io_in_4_bits_payload_g_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( T16 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_g_type( io_in_3_bits_payload_g_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T14 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T12 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T10 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_3_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_3_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_3_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_3_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_g_type( LockingRRArbiter_3_io_out_bits_payload_g_type ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_8 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_4_io_in_4_ready ),
       .io_in_4_valid( T8 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_addr_beat( io_in_4_bits_payload_addr_beat ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_is_builtin_type( io_in_4_bits_payload_is_builtin_type ),
       .io_in_4_bits_payload_g_type( io_in_4_bits_payload_g_type ),
       .io_in_4_bits_payload_data( io_in_4_bits_payload_data ),
       .io_in_3_ready( LockingRRArbiter_4_io_in_3_ready ),
       .io_in_3_valid( T6 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_addr_beat( io_in_3_bits_payload_addr_beat ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_is_builtin_type( io_in_3_bits_payload_is_builtin_type ),
       .io_in_3_bits_payload_g_type( io_in_3_bits_payload_g_type ),
       .io_in_3_bits_payload_data( io_in_3_bits_payload_data ),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( io_in_2_bits_payload_addr_beat ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_is_builtin_type( io_in_2_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( io_in_1_bits_payload_addr_beat ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_is_builtin_type( io_in_1_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( io_in_0_bits_payload_addr_beat ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_is_builtin_type( io_in_0_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_out_ready( io_out_4_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_4_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_4_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_4_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_g_type( LockingRRArbiter_4_io_out_bits_payload_g_type ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_9(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [3:0] io_in_4_bits_payload_manager_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [3:0] io_in_3_bits_payload_manager_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_header_src,
    output[2:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire T7;
  wire T8;
  reg [2:0] last_grant;
  wire[2:0] T124;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire T20;
  wire[2:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T15 ? 3'h1 : T0;
  assign T0 = T13 ? 3'h2 : T1;
  assign T1 = T11 ? 3'h3 : T2;
  assign T2 = T7 ? 3'h4 : T3;
  assign T3 = io_in_0_valid ? 3'h0 : T4;
  assign T4 = io_in_1_valid ? 3'h1 : T5;
  assign T5 = io_in_2_valid ? 3'h2 : T6;
  assign T6 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T7 = io_in_4_valid & T8;
  assign T8 = last_grant < 3'h4;
  assign T124 = reset ? 3'h0 : T9;
  assign T9 = T10 ? chosen : last_grant;
  assign T10 = io_out_ready & io_out_valid;
  assign T11 = io_in_3_valid & T12;
  assign T12 = last_grant < 3'h3;
  assign T13 = io_in_2_valid & T14;
  assign T14 = last_grant < 3'h2;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 3'h1;
  assign io_out_bits_payload_manager_xact_id = T17;
  assign T17 = T25 ? io_in_4_bits_payload_manager_xact_id : T18;
  assign T18 = T24 ? T22 : T19;
  assign T19 = T20 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T20 = T21[1'h0];
  assign T21 = chosen;
  assign T22 = T23 ? io_in_3_bits_payload_manager_xact_id : io_in_2_bits_payload_manager_xact_id;
  assign T23 = T21[1'h0];
  assign T24 = T21[1'h1];
  assign T25 = T21[2'h2];
  assign io_out_bits_header_dst = T26;
  assign T26 = T33 ? io_in_4_bits_header_dst : T27;
  assign T27 = T32 ? T30 : T28;
  assign T28 = T29 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T29 = T21[1'h0];
  assign T30 = T31 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T31 = T21[1'h0];
  assign T32 = T21[1'h1];
  assign T33 = T21[2'h2];
  assign io_out_bits_header_src = T34;
  assign T34 = T41 ? io_in_4_bits_header_src : T35;
  assign T35 = T40 ? T38 : T36;
  assign T36 = T37 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T37 = T21[1'h0];
  assign T38 = T39 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T39 = T21[1'h0];
  assign T40 = T21[1'h1];
  assign T41 = T21[2'h2];
  assign io_out_valid = T42;
  assign T42 = T49 ? io_in_4_valid : T43;
  assign T43 = T48 ? T46 : T44;
  assign T44 = T45 ? io_in_1_valid : io_in_0_valid;
  assign T45 = T21[1'h0];
  assign T46 = T47 ? io_in_3_valid : io_in_2_valid;
  assign T47 = T21[1'h0];
  assign T48 = T21[1'h1];
  assign T49 = T21[2'h2];
  assign io_in_0_ready = T50;
  assign T50 = T51 & io_out_ready;
  assign T51 = T67 | T52;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T56 | T54;
  assign T54 = io_in_4_valid & T55;
  assign T55 = last_grant < 3'h4;
  assign T56 = T59 | T57;
  assign T57 = io_in_3_valid & T58;
  assign T58 = last_grant < 3'h3;
  assign T59 = T62 | T60;
  assign T60 = io_in_2_valid & T61;
  assign T61 = last_grant < 3'h2;
  assign T62 = T65 | T63;
  assign T63 = io_in_1_valid & T64;
  assign T64 = last_grant < 3'h1;
  assign T65 = io_in_0_valid & T66;
  assign T66 = last_grant < 3'h0;
  assign T67 = last_grant < 3'h0;
  assign io_in_1_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = T76 | T70;
  assign T70 = T71 ^ 1'h1;
  assign T71 = T72 | io_in_0_valid;
  assign T72 = T73 | T54;
  assign T73 = T74 | T57;
  assign T74 = T75 | T60;
  assign T75 = T65 | T63;
  assign T76 = T78 & T77;
  assign T77 = last_grant < 3'h1;
  assign T78 = T65 ^ 1'h1;
  assign io_in_2_ready = T79;
  assign T79 = T80 & io_out_ready;
  assign T80 = T88 | T81;
  assign T81 = T82 ^ 1'h1;
  assign T82 = T83 | io_in_1_valid;
  assign T83 = T84 | io_in_0_valid;
  assign T84 = T85 | T54;
  assign T85 = T86 | T57;
  assign T86 = T87 | T60;
  assign T87 = T65 | T63;
  assign T88 = T90 & T89;
  assign T89 = last_grant < 3'h2;
  assign T90 = T91 ^ 1'h1;
  assign T91 = T65 | T63;
  assign io_in_3_ready = T92;
  assign T92 = T93 & io_out_ready;
  assign T93 = T102 | T94;
  assign T94 = T95 ^ 1'h1;
  assign T95 = T96 | io_in_2_valid;
  assign T96 = T97 | io_in_1_valid;
  assign T97 = T98 | io_in_0_valid;
  assign T98 = T99 | T54;
  assign T99 = T100 | T57;
  assign T100 = T101 | T60;
  assign T101 = T65 | T63;
  assign T102 = T104 & T103;
  assign T103 = last_grant < 3'h3;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T106 | T60;
  assign T106 = T65 | T63;
  assign io_in_4_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = T118 | T109;
  assign T109 = T110 ^ 1'h1;
  assign T110 = T111 | io_in_3_valid;
  assign T111 = T112 | io_in_2_valid;
  assign T112 = T113 | io_in_1_valid;
  assign T113 = T114 | io_in_0_valid;
  assign T114 = T115 | T54;
  assign T115 = T116 | T57;
  assign T116 = T117 | T60;
  assign T117 = T65 | T63;
  assign T118 = T120 & T119;
  assign T119 = last_grant < 3'h4;
  assign T120 = T121 ^ 1'h1;
  assign T121 = T122 | T57;
  assign T122 = T123 | T60;
  assign T123 = T65 | T63;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T10) begin
      last_grant <= chosen;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [2:0] io_in_4_bits_header_src,
    input [2:0] io_in_4_bits_header_dst,
    input [3:0] io_in_4_bits_payload_manager_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [2:0] io_in_3_bits_header_src,
    input [2:0] io_in_3_bits_header_dst,
    input [3:0] io_in_3_bits_payload_manager_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [2:0] io_in_2_bits_header_src,
    input [2:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_header_src,
    input [2:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_header_src,
    input [2:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_4_ready,
    output io_out_4_valid,
    output[2:0] io_out_4_bits_header_src,
    output[2:0] io_out_4_bits_header_dst,
    output[3:0] io_out_4_bits_payload_manager_xact_id,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[2:0] io_out_3_bits_header_src,
    output[2:0] io_out_3_bits_header_dst,
    output[3:0] io_out_3_bits_payload_manager_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[2:0] io_out_2_bits_header_src,
    output[2:0] io_out_2_bits_header_dst,
    output[3:0] io_out_2_bits_payload_manager_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[2:0] io_out_1_bits_header_src,
    output[2:0] io_out_1_bits_header_dst,
    output[3:0] io_out_1_bits_payload_manager_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[2:0] io_out_0_bits_header_src,
    output[2:0] io_out_0_bits_header_dst,
    output[3:0] io_out_0_bits_payload_manager_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[2:0] LockingRRArbiter_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_2_io_in_4_ready;
  wire LockingRRArbiter_2_io_in_3_ready;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_3_io_in_4_ready;
  wire LockingRRArbiter_3_io_in_3_ready;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_3_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_4_io_in_4_ready;
  wire LockingRRArbiter_4_io_in_3_ready;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[2:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_4_io_out_bits_payload_manager_xact_id;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 3'h4;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 3'h4;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 3'h4;
  assign T6 = io_in_3_valid & T7;
  assign T7 = io_in_3_bits_header_dst == 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = io_in_4_bits_header_dst == 3'h4;
  assign T10 = io_in_0_valid & T11;
  assign T11 = io_in_0_bits_header_dst == 3'h3;
  assign T12 = io_in_1_valid & T13;
  assign T13 = io_in_1_bits_header_dst == 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = io_in_2_bits_header_dst == 3'h3;
  assign T16 = io_in_3_valid & T17;
  assign T17 = io_in_3_bits_header_dst == 3'h3;
  assign T18 = io_in_4_valid & T19;
  assign T19 = io_in_4_bits_header_dst == 3'h3;
  assign T20 = io_in_0_valid & T21;
  assign T21 = io_in_0_bits_header_dst == 3'h2;
  assign T22 = io_in_1_valid & T23;
  assign T23 = io_in_1_bits_header_dst == 3'h2;
  assign T24 = io_in_2_valid & T25;
  assign T25 = io_in_2_bits_header_dst == 3'h2;
  assign T26 = io_in_3_valid & T27;
  assign T27 = io_in_3_bits_header_dst == 3'h2;
  assign T28 = io_in_4_valid & T29;
  assign T29 = io_in_4_bits_header_dst == 3'h2;
  assign T30 = io_in_0_valid & T31;
  assign T31 = io_in_0_bits_header_dst == 3'h1;
  assign T32 = io_in_1_valid & T33;
  assign T33 = io_in_1_bits_header_dst == 3'h1;
  assign T34 = io_in_2_valid & T35;
  assign T35 = io_in_2_bits_header_dst == 3'h1;
  assign T36 = io_in_3_valid & T37;
  assign T37 = io_in_3_bits_header_dst == 3'h1;
  assign T38 = io_in_4_valid & T39;
  assign T39 = io_in_4_bits_header_dst == 3'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = io_in_0_bits_header_dst == 3'h0;
  assign T42 = io_in_1_valid & T43;
  assign T43 = io_in_1_bits_header_dst == 3'h0;
  assign T44 = io_in_2_valid & T45;
  assign T45 = io_in_2_bits_header_dst == 3'h0;
  assign T46 = io_in_3_valid & T47;
  assign T47 = io_in_3_bits_header_dst == 3'h0;
  assign T48 = io_in_4_valid & T49;
  assign T49 = io_in_4_bits_header_dst == 3'h0;
  assign io_out_0_bits_payload_manager_xact_id = LockingRRArbiter_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_io_out_valid;
  assign io_out_1_bits_payload_manager_xact_id = LockingRRArbiter_1_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_manager_xact_id = LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_out_3_bits_payload_manager_xact_id = LockingRRArbiter_3_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_3_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_3_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_4_bits_payload_manager_xact_id = LockingRRArbiter_4_io_out_bits_payload_manager_xact_id;
  assign io_out_4_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_4_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_4_valid = LockingRRArbiter_4_io_out_valid;
  assign io_in_0_ready = T50;
  assign T50 = T54 | T51;
  assign T51 = T52;
  assign T52 = LockingRRArbiter_4_io_in_0_ready & T53;
  assign T53 = io_in_0_bits_header_dst == 3'h4;
  assign T54 = T58 | T55;
  assign T55 = T56;
  assign T56 = LockingRRArbiter_3_io_in_0_ready & T57;
  assign T57 = io_in_0_bits_header_dst == 3'h3;
  assign T58 = T62 | T59;
  assign T59 = T60;
  assign T60 = LockingRRArbiter_2_io_in_0_ready & T61;
  assign T61 = io_in_0_bits_header_dst == 3'h2;
  assign T62 = T66 | T63;
  assign T63 = T64;
  assign T64 = LockingRRArbiter_1_io_in_0_ready & T65;
  assign T65 = io_in_0_bits_header_dst == 3'h1;
  assign T66 = T67;
  assign T67 = LockingRRArbiter_io_in_0_ready & T68;
  assign T68 = io_in_0_bits_header_dst == 3'h0;
  assign io_in_1_ready = T69;
  assign T69 = T73 | T70;
  assign T70 = T71;
  assign T71 = LockingRRArbiter_4_io_in_1_ready & T72;
  assign T72 = io_in_1_bits_header_dst == 3'h4;
  assign T73 = T77 | T74;
  assign T74 = T75;
  assign T75 = LockingRRArbiter_3_io_in_1_ready & T76;
  assign T76 = io_in_1_bits_header_dst == 3'h3;
  assign T77 = T81 | T78;
  assign T78 = T79;
  assign T79 = LockingRRArbiter_2_io_in_1_ready & T80;
  assign T80 = io_in_1_bits_header_dst == 3'h2;
  assign T81 = T85 | T82;
  assign T82 = T83;
  assign T83 = LockingRRArbiter_1_io_in_1_ready & T84;
  assign T84 = io_in_1_bits_header_dst == 3'h1;
  assign T85 = T86;
  assign T86 = LockingRRArbiter_io_in_1_ready & T87;
  assign T87 = io_in_1_bits_header_dst == 3'h0;
  assign io_in_2_ready = T88;
  assign T88 = T92 | T89;
  assign T89 = T90;
  assign T90 = LockingRRArbiter_4_io_in_2_ready & T91;
  assign T91 = io_in_2_bits_header_dst == 3'h4;
  assign T92 = T96 | T93;
  assign T93 = T94;
  assign T94 = LockingRRArbiter_3_io_in_2_ready & T95;
  assign T95 = io_in_2_bits_header_dst == 3'h3;
  assign T96 = T100 | T97;
  assign T97 = T98;
  assign T98 = LockingRRArbiter_2_io_in_2_ready & T99;
  assign T99 = io_in_2_bits_header_dst == 3'h2;
  assign T100 = T104 | T101;
  assign T101 = T102;
  assign T102 = LockingRRArbiter_1_io_in_2_ready & T103;
  assign T103 = io_in_2_bits_header_dst == 3'h1;
  assign T104 = T105;
  assign T105 = LockingRRArbiter_io_in_2_ready & T106;
  assign T106 = io_in_2_bits_header_dst == 3'h0;
  assign io_in_3_ready = T107;
  assign T107 = T111 | T108;
  assign T108 = T109;
  assign T109 = LockingRRArbiter_4_io_in_3_ready & T110;
  assign T110 = io_in_3_bits_header_dst == 3'h4;
  assign T111 = T115 | T112;
  assign T112 = T113;
  assign T113 = LockingRRArbiter_3_io_in_3_ready & T114;
  assign T114 = io_in_3_bits_header_dst == 3'h3;
  assign T115 = T119 | T116;
  assign T116 = T117;
  assign T117 = LockingRRArbiter_2_io_in_3_ready & T118;
  assign T118 = io_in_3_bits_header_dst == 3'h2;
  assign T119 = T123 | T120;
  assign T120 = T121;
  assign T121 = LockingRRArbiter_1_io_in_3_ready & T122;
  assign T122 = io_in_3_bits_header_dst == 3'h1;
  assign T123 = T124;
  assign T124 = LockingRRArbiter_io_in_3_ready & T125;
  assign T125 = io_in_3_bits_header_dst == 3'h0;
  assign io_in_4_ready = T126;
  assign T126 = T130 | T127;
  assign T127 = T128;
  assign T128 = LockingRRArbiter_4_io_in_4_ready & T129;
  assign T129 = io_in_4_bits_header_dst == 3'h4;
  assign T130 = T134 | T131;
  assign T131 = T132;
  assign T132 = LockingRRArbiter_3_io_in_4_ready & T133;
  assign T133 = io_in_4_bits_header_dst == 3'h3;
  assign T134 = T138 | T135;
  assign T135 = T136;
  assign T136 = LockingRRArbiter_2_io_in_4_ready & T137;
  assign T137 = io_in_4_bits_header_dst == 3'h2;
  assign T138 = T142 | T139;
  assign T139 = T140;
  assign T140 = LockingRRArbiter_1_io_in_4_ready & T141;
  assign T141 = io_in_4_bits_header_dst == 3'h1;
  assign T142 = T143;
  assign T143 = LockingRRArbiter_io_in_4_ready & T144;
  assign T144 = io_in_4_bits_header_dst == 3'h0;
  LockingRRArbiter_9 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( T48 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( T46 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( T44 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( T42 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( T38 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( T36 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T34 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T32 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T30 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_1_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( T28 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_3_ready( LockingRRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( T26 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T24 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T22 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_2_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( T18 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_3_ready( LockingRRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( T16 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T14 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T12 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T10 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_3_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_3_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_4_io_in_4_ready ),
       .io_in_4_valid( T8 ),
       .io_in_4_bits_header_src( io_in_4_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_bits_payload_manager_xact_id ),
       .io_in_3_ready( LockingRRArbiter_4_io_in_3_ready ),
       .io_in_3_valid( T6 ),
       .io_in_3_bits_header_src( io_in_3_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_bits_payload_manager_xact_id ),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_4_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_4_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipTileLinkCrossbar(input clk, input reset,
    output io_clients_2_acquire_ready,
    input  io_clients_2_acquire_valid,
    input [25:0] io_clients_2_acquire_bits_addr_block,
    input [5:0] io_clients_2_acquire_bits_client_xact_id,
    input [1:0] io_clients_2_acquire_bits_addr_beat,
    input  io_clients_2_acquire_bits_is_builtin_type,
    input [2:0] io_clients_2_acquire_bits_a_type,
    input [16:0] io_clients_2_acquire_bits_union,
    input [127:0] io_clients_2_acquire_bits_data,
    input  io_clients_2_grant_ready,
    output io_clients_2_grant_valid,
    output[1:0] io_clients_2_grant_bits_addr_beat,
    output[5:0] io_clients_2_grant_bits_client_xact_id,
    output[3:0] io_clients_2_grant_bits_manager_xact_id,
    output io_clients_2_grant_bits_is_builtin_type,
    output[3:0] io_clients_2_grant_bits_g_type,
    output[127:0] io_clients_2_grant_bits_data,
    input  io_clients_2_probe_ready,
    output io_clients_2_probe_valid,
    output[25:0] io_clients_2_probe_bits_addr_block,
    output[1:0] io_clients_2_probe_bits_p_type,
    output io_clients_2_release_ready,
    input  io_clients_2_release_valid,
    input [1:0] io_clients_2_release_bits_addr_beat,
    input [25:0] io_clients_2_release_bits_addr_block,
    input [5:0] io_clients_2_release_bits_client_xact_id,
    input  io_clients_2_release_bits_voluntary,
    input [2:0] io_clients_2_release_bits_r_type,
    input [127:0] io_clients_2_release_bits_data,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [25:0] io_clients_1_acquire_bits_addr_block,
    input [5:0] io_clients_1_acquire_bits_client_xact_id,
    input [1:0] io_clients_1_acquire_bits_addr_beat,
    input  io_clients_1_acquire_bits_is_builtin_type,
    input [2:0] io_clients_1_acquire_bits_a_type,
    input [16:0] io_clients_1_acquire_bits_union,
    input [127:0] io_clients_1_acquire_bits_data,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_addr_beat,
    output[5:0] io_clients_1_grant_bits_client_xact_id,
    output[3:0] io_clients_1_grant_bits_manager_xact_id,
    output io_clients_1_grant_bits_is_builtin_type,
    output[3:0] io_clients_1_grant_bits_g_type,
    output[127:0] io_clients_1_grant_bits_data,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[25:0] io_clients_1_probe_bits_addr_block,
    output[1:0] io_clients_1_probe_bits_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_addr_beat,
    input [25:0] io_clients_1_release_bits_addr_block,
    input [5:0] io_clients_1_release_bits_client_xact_id,
    input  io_clients_1_release_bits_voluntary,
    input [2:0] io_clients_1_release_bits_r_type,
    input [127:0] io_clients_1_release_bits_data,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [25:0] io_clients_0_acquire_bits_addr_block,
    input [5:0] io_clients_0_acquire_bits_client_xact_id,
    input [1:0] io_clients_0_acquire_bits_addr_beat,
    input  io_clients_0_acquire_bits_is_builtin_type,
    input [2:0] io_clients_0_acquire_bits_a_type,
    input [16:0] io_clients_0_acquire_bits_union,
    input [127:0] io_clients_0_acquire_bits_data,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_addr_beat,
    output[5:0] io_clients_0_grant_bits_client_xact_id,
    output[3:0] io_clients_0_grant_bits_manager_xact_id,
    output io_clients_0_grant_bits_is_builtin_type,
    output[3:0] io_clients_0_grant_bits_g_type,
    output[127:0] io_clients_0_grant_bits_data,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[25:0] io_clients_0_probe_bits_addr_block,
    output[1:0] io_clients_0_probe_bits_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_addr_beat,
    input [25:0] io_clients_0_release_bits_addr_block,
    input [5:0] io_clients_0_release_bits_client_xact_id,
    input  io_clients_0_release_bits_voluntary,
    input [2:0] io_clients_0_release_bits_r_type,
    input [127:0] io_clients_0_release_bits_data,
    input  io_managers_1_acquire_ready,
    output io_managers_1_acquire_valid,
    output[25:0] io_managers_1_acquire_bits_addr_block,
    output[5:0] io_managers_1_acquire_bits_client_xact_id,
    output[1:0] io_managers_1_acquire_bits_addr_beat,
    output io_managers_1_acquire_bits_is_builtin_type,
    output[2:0] io_managers_1_acquire_bits_a_type,
    output[16:0] io_managers_1_acquire_bits_union,
    output[127:0] io_managers_1_acquire_bits_data,
    output[1:0] io_managers_1_acquire_bits_client_id,
    output io_managers_1_grant_ready,
    input  io_managers_1_grant_valid,
    input [1:0] io_managers_1_grant_bits_addr_beat,
    input [5:0] io_managers_1_grant_bits_client_xact_id,
    input [3:0] io_managers_1_grant_bits_manager_xact_id,
    input  io_managers_1_grant_bits_is_builtin_type,
    input [3:0] io_managers_1_grant_bits_g_type,
    input [127:0] io_managers_1_grant_bits_data,
    input [1:0] io_managers_1_grant_bits_client_id,
    input  io_managers_1_finish_ready,
    output io_managers_1_finish_valid,
    output[3:0] io_managers_1_finish_bits_manager_xact_id,
    output io_managers_1_probe_ready,
    input  io_managers_1_probe_valid,
    input [25:0] io_managers_1_probe_bits_addr_block,
    input [1:0] io_managers_1_probe_bits_p_type,
    input [1:0] io_managers_1_probe_bits_client_id,
    input  io_managers_1_release_ready,
    output io_managers_1_release_valid,
    output[1:0] io_managers_1_release_bits_addr_beat,
    output[25:0] io_managers_1_release_bits_addr_block,
    output[5:0] io_managers_1_release_bits_client_xact_id,
    output io_managers_1_release_bits_voluntary,
    output[2:0] io_managers_1_release_bits_r_type,
    output[127:0] io_managers_1_release_bits_data,
    output[1:0] io_managers_1_release_bits_client_id,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[25:0] io_managers_0_acquire_bits_addr_block,
    output[5:0] io_managers_0_acquire_bits_client_xact_id,
    output[1:0] io_managers_0_acquire_bits_addr_beat,
    output io_managers_0_acquire_bits_is_builtin_type,
    output[2:0] io_managers_0_acquire_bits_a_type,
    output[16:0] io_managers_0_acquire_bits_union,
    output[127:0] io_managers_0_acquire_bits_data,
    output[1:0] io_managers_0_acquire_bits_client_id,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_addr_beat,
    input [5:0] io_managers_0_grant_bits_client_xact_id,
    input [3:0] io_managers_0_grant_bits_manager_xact_id,
    input  io_managers_0_grant_bits_is_builtin_type,
    input [3:0] io_managers_0_grant_bits_g_type,
    input [127:0] io_managers_0_grant_bits_data,
    input [1:0] io_managers_0_grant_bits_client_id,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output[3:0] io_managers_0_finish_bits_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [25:0] io_managers_0_probe_bits_addr_block,
    input [1:0] io_managers_0_probe_bits_p_type,
    input [1:0] io_managers_0_probe_bits_client_id,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[1:0] io_managers_0_release_bits_addr_beat,
    output[25:0] io_managers_0_release_bits_addr_block,
    output[5:0] io_managers_0_release_bits_client_xact_id,
    output io_managers_0_release_bits_voluntary,
    output[2:0] io_managers_0_release_bits_r_type,
    output[127:0] io_managers_0_release_bits_data,
    output[1:0] io_managers_0_release_bits_client_id
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire T6;
  wire[3:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[3:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[127:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[3:0] T23;
  wire[5:0] T24;
  wire[1:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire T29;
  wire[127:0] T30;
  wire[3:0] T31;
  wire T32;
  wire[3:0] T33;
  wire[5:0] T34;
  wire[1:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[1:0] T43;
  wire[25:0] T44;
  wire[2:0] T45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire T48;
  wire[1:0] T49;
  wire[25:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[127:0] T57;
  wire[2:0] T58;
  wire T59;
  wire[5:0] T60;
  wire[25:0] T61;
  wire[1:0] T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire[2:0] T65;
  wire T66;
  wire[127:0] T67;
  wire[2:0] T68;
  wire T69;
  wire[5:0] T70;
  wire[25:0] T71;
  wire[1:0] T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire T76;
  wire[127:0] T77;
  wire[2:0] T78;
  wire T79;
  wire[5:0] T80;
  wire[25:0] T81;
  wire[1:0] T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[127:0] T89;
  wire[16:0] T90;
  wire[2:0] T91;
  wire T92;
  wire[1:0] T93;
  wire[5:0] T94;
  wire[25:0] T95;
  wire[2:0] T96;
  wire[2:0] T97;
  wire[2:0] T98;
  wire T99;
  wire[127:0] T100;
  wire[16:0] T101;
  wire[2:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[5:0] T105;
  wire[25:0] T106;
  wire[2:0] T107;
  wire[2:0] T108;
  wire[2:0] T109;
  wire T110;
  wire[127:0] T111;
  wire[16:0] T112;
  wire[2:0] T113;
  wire T114;
  wire[1:0] T115;
  wire[5:0] T116;
  wire[25:0] T117;
  wire[2:0] T118;
  wire[2:0] T119;
  wire[2:0] T120;
  wire T121;
  wire[127:0] T122;
  wire[2:0] T123;
  wire T124;
  wire[5:0] T125;
  wire[25:0] T126;
  wire[1:0] T127;
  wire[2:0] T128;
  wire[2:0] T129;
  wire[2:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[2:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  wire T138;
  wire[127:0] T139;
  wire[16:0] T140;
  wire[2:0] T141;
  wire T142;
  wire[1:0] T143;
  wire[5:0] T144;
  wire[25:0] T145;
  wire[2:0] T146;
  wire[2:0] T147;
  wire[2:0] T148;
  wire T149;
  wire[127:0] T150;
  wire[2:0] T151;
  wire T152;
  wire[5:0] T153;
  wire[25:0] T154;
  wire[1:0] T155;
  wire[2:0] T156;
  wire[2:0] T157;
  wire[2:0] T158;
  wire T159;
  wire T160;
  wire[3:0] T161;
  wire[2:0] T162;
  wire[2:0] T163;
  wire[2:0] T164;
  wire T165;
  wire T166;
  wire[127:0] T167;
  wire[16:0] T168;
  wire[2:0] T169;
  wire T170;
  wire[1:0] T171;
  wire[5:0] T172;
  wire[25:0] T173;
  wire[2:0] T174;
  wire[2:0] T175;
  wire[2:0] T176;
  wire T177;
  wire T178;
  wire[1:0] T179;
  wire[25:0] T180;
  wire[2:0] T181;
  wire[2:0] T182;
  wire[2:0] T183;
  wire T184;
  wire T185;
  wire[127:0] T186;
  wire[3:0] T187;
  wire T188;
  wire[3:0] T189;
  wire[5:0] T190;
  wire[1:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire[1:0] T198;
  wire[25:0] T199;
  wire[2:0] T200;
  wire[2:0] T201;
  wire[2:0] T202;
  wire T203;
  wire T204;
  wire[127:0] T205;
  wire[3:0] T206;
  wire T207;
  wire[3:0] T208;
  wire[5:0] T209;
  wire[1:0] T210;
  wire[2:0] T211;
  wire[2:0] T212;
  wire[2:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[1:0] T217;
  wire[25:0] T218;
  wire[2:0] T219;
  wire[2:0] T220;
  wire[2:0] T221;
  wire T222;
  wire T223;
  wire[127:0] T224;
  wire[3:0] T225;
  wire T226;
  wire[3:0] T227;
  wire[5:0] T228;
  wire[1:0] T229;
  wire[2:0] T230;
  wire[2:0] T231;
  wire[2:0] T232;
  wire T233;
  wire T234;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  wire[5:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_io_manager_finish_valid;
  wire[3:0] ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_io_manager_release_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  wire[5:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_io_network_grant_valid;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_src;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat;
  wire[5:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type;
  wire[127:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data;
  wire ManagerTileLinkNetworkPort_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_io_network_probe_valid;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_src;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_io_network_release_ready;
  wire ManagerTileLinkNetworkPort_1_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_block;
  wire[5:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_beat;
  wire ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_union;
  wire[127:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_1_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_1_io_manager_finish_valid;
  wire[3:0] ManagerTileLinkNetworkPort_1_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_1_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_1_io_manager_release_valid;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_beat;
  wire[25:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_block;
  wire[5:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_xact_id;
  wire ManagerTileLinkNetworkPort_1_io_manager_release_bits_voluntary;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_r_type;
  wire[127:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_1_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_1_io_network_grant_valid;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire[5:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire[3:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire[127:0] ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire ManagerTileLinkNetworkPort_1_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_1_io_network_probe_valid;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire[2:0] ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_1_io_network_release_ready;
  wire TileLinkEnqueuer_io_client_acquire_ready;
  wire TileLinkEnqueuer_io_client_grant_valid;
  wire[2:0] TileLinkEnqueuer_io_client_grant_bits_header_src;
  wire[2:0] TileLinkEnqueuer_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat;
  wire[5:0] TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_io_client_finish_ready;
  wire TileLinkEnqueuer_io_client_probe_valid;
  wire[2:0] TileLinkEnqueuer_io_client_probe_bits_header_src;
  wire[2:0] TileLinkEnqueuer_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_io_client_release_ready;
  wire TileLinkEnqueuer_io_manager_acquire_valid;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_header_src;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_io_manager_grant_ready;
  wire TileLinkEnqueuer_io_manager_finish_valid;
  wire[2:0] TileLinkEnqueuer_io_manager_finish_bits_header_src;
  wire[2:0] TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_manager_probe_ready;
  wire TileLinkEnqueuer_io_manager_release_valid;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_header_src;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_acquire_ready;
  wire TileLinkEnqueuer_1_io_client_grant_valid;
  wire[2:0] TileLinkEnqueuer_1_io_client_grant_bits_header_src;
  wire[2:0] TileLinkEnqueuer_1_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat;
  wire[5:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_finish_ready;
  wire TileLinkEnqueuer_1_io_client_probe_valid;
  wire[2:0] TileLinkEnqueuer_1_io_client_probe_bits_header_src;
  wire[2:0] TileLinkEnqueuer_1_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_1_io_client_release_ready;
  wire TileLinkEnqueuer_1_io_manager_acquire_valid;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_src;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_1_io_manager_grant_ready;
  wire TileLinkEnqueuer_1_io_manager_finish_valid;
  wire[2:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_src;
  wire[2:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_manager_probe_ready;
  wire TileLinkEnqueuer_1_io_manager_release_valid;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_header_src;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_acquire_ready;
  wire TileLinkEnqueuer_2_io_client_grant_valid;
  wire[2:0] TileLinkEnqueuer_2_io_client_grant_bits_header_src;
  wire[2:0] TileLinkEnqueuer_2_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat;
  wire[5:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_finish_ready;
  wire TileLinkEnqueuer_2_io_client_probe_valid;
  wire[2:0] TileLinkEnqueuer_2_io_client_probe_bits_header_src;
  wire[2:0] TileLinkEnqueuer_2_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_2_io_client_release_ready;
  wire TileLinkEnqueuer_2_io_manager_acquire_valid;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_src;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_2_io_manager_grant_ready;
  wire TileLinkEnqueuer_2_io_manager_finish_valid;
  wire[2:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_src;
  wire[2:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_manager_probe_ready;
  wire TileLinkEnqueuer_2_io_manager_release_valid;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_header_src;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_acquire_ready;
  wire TileLinkEnqueuer_3_io_client_grant_valid;
  wire[2:0] TileLinkEnqueuer_3_io_client_grant_bits_header_src;
  wire[2:0] TileLinkEnqueuer_3_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat;
  wire[5:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_finish_ready;
  wire TileLinkEnqueuer_3_io_client_probe_valid;
  wire[2:0] TileLinkEnqueuer_3_io_client_probe_bits_header_src;
  wire[2:0] TileLinkEnqueuer_3_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_3_io_client_release_ready;
  wire TileLinkEnqueuer_3_io_manager_acquire_valid;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_src;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_3_io_manager_grant_ready;
  wire TileLinkEnqueuer_3_io_manager_finish_valid;
  wire[2:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_src;
  wire[2:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_manager_probe_ready;
  wire TileLinkEnqueuer_3_io_manager_release_valid;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_header_src;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_4_io_client_acquire_ready;
  wire TileLinkEnqueuer_4_io_client_grant_valid;
  wire[2:0] TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  wire[2:0] TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  wire[5:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_4_io_client_finish_ready;
  wire TileLinkEnqueuer_4_io_client_probe_valid;
  wire[2:0] TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  wire[2:0] TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_4_io_client_release_ready;
  wire TileLinkEnqueuer_4_io_manager_acquire_valid;
  wire[2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_src;
  wire[2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_4_io_manager_grant_ready;
  wire TileLinkEnqueuer_4_io_manager_finish_valid;
  wire[2:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_src;
  wire[2:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  wire[3:0] TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_4_io_manager_probe_ready;
  wire TileLinkEnqueuer_4_io_manager_release_valid;
  wire[2:0] TileLinkEnqueuer_4_io_manager_release_bits_header_src;
  wire[2:0] TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  wire[5:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  wire acqNet_io_in_4_ready;
  wire acqNet_io_in_3_ready;
  wire acqNet_io_in_2_ready;
  wire acqNet_io_out_1_valid;
  wire[2:0] acqNet_io_out_1_bits_header_src;
  wire[2:0] acqNet_io_out_1_bits_header_dst;
  wire[25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire[5:0] acqNet_io_out_1_bits_payload_client_xact_id;
  wire[1:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire acqNet_io_out_1_bits_payload_is_builtin_type;
  wire[2:0] acqNet_io_out_1_bits_payload_a_type;
  wire[16:0] acqNet_io_out_1_bits_payload_union;
  wire[127:0] acqNet_io_out_1_bits_payload_data;
  wire acqNet_io_out_0_valid;
  wire[2:0] acqNet_io_out_0_bits_header_src;
  wire[2:0] acqNet_io_out_0_bits_header_dst;
  wire[25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire[5:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[1:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire acqNet_io_out_0_bits_payload_is_builtin_type;
  wire[2:0] acqNet_io_out_0_bits_payload_a_type;
  wire[16:0] acqNet_io_out_0_bits_payload_union;
  wire[127:0] acqNet_io_out_0_bits_payload_data;
  wire relNet_io_in_4_ready;
  wire relNet_io_in_3_ready;
  wire relNet_io_in_2_ready;
  wire relNet_io_out_1_valid;
  wire[2:0] relNet_io_out_1_bits_header_src;
  wire[2:0] relNet_io_out_1_bits_header_dst;
  wire[1:0] relNet_io_out_1_bits_payload_addr_beat;
  wire[25:0] relNet_io_out_1_bits_payload_addr_block;
  wire[5:0] relNet_io_out_1_bits_payload_client_xact_id;
  wire relNet_io_out_1_bits_payload_voluntary;
  wire[2:0] relNet_io_out_1_bits_payload_r_type;
  wire[127:0] relNet_io_out_1_bits_payload_data;
  wire relNet_io_out_0_valid;
  wire[2:0] relNet_io_out_0_bits_header_src;
  wire[2:0] relNet_io_out_0_bits_header_dst;
  wire[1:0] relNet_io_out_0_bits_payload_addr_beat;
  wire[25:0] relNet_io_out_0_bits_payload_addr_block;
  wire[5:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire relNet_io_out_0_bits_payload_voluntary;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire[127:0] relNet_io_out_0_bits_payload_data;
  wire prbNet_io_in_1_ready;
  wire prbNet_io_in_0_ready;
  wire prbNet_io_out_4_valid;
  wire[2:0] prbNet_io_out_4_bits_header_src;
  wire[2:0] prbNet_io_out_4_bits_header_dst;
  wire[25:0] prbNet_io_out_4_bits_payload_addr_block;
  wire[1:0] prbNet_io_out_4_bits_payload_p_type;
  wire prbNet_io_out_3_valid;
  wire[2:0] prbNet_io_out_3_bits_header_src;
  wire[2:0] prbNet_io_out_3_bits_header_dst;
  wire[25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire[1:0] prbNet_io_out_3_bits_payload_p_type;
  wire prbNet_io_out_2_valid;
  wire[2:0] prbNet_io_out_2_bits_header_src;
  wire[2:0] prbNet_io_out_2_bits_header_dst;
  wire[25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire gntNet_io_in_1_ready;
  wire gntNet_io_in_0_ready;
  wire gntNet_io_out_4_valid;
  wire[2:0] gntNet_io_out_4_bits_header_src;
  wire[2:0] gntNet_io_out_4_bits_header_dst;
  wire[1:0] gntNet_io_out_4_bits_payload_addr_beat;
  wire[5:0] gntNet_io_out_4_bits_payload_client_xact_id;
  wire[3:0] gntNet_io_out_4_bits_payload_manager_xact_id;
  wire gntNet_io_out_4_bits_payload_is_builtin_type;
  wire[3:0] gntNet_io_out_4_bits_payload_g_type;
  wire[127:0] gntNet_io_out_4_bits_payload_data;
  wire gntNet_io_out_3_valid;
  wire[2:0] gntNet_io_out_3_bits_header_src;
  wire[2:0] gntNet_io_out_3_bits_header_dst;
  wire[1:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire[5:0] gntNet_io_out_3_bits_payload_client_xact_id;
  wire[3:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire gntNet_io_out_3_bits_payload_is_builtin_type;
  wire[3:0] gntNet_io_out_3_bits_payload_g_type;
  wire[127:0] gntNet_io_out_3_bits_payload_data;
  wire gntNet_io_out_2_valid;
  wire[2:0] gntNet_io_out_2_bits_header_src;
  wire[2:0] gntNet_io_out_2_bits_header_dst;
  wire[1:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire[5:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[3:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire gntNet_io_out_2_bits_payload_is_builtin_type;
  wire[3:0] gntNet_io_out_2_bits_payload_g_type;
  wire[127:0] gntNet_io_out_2_bits_payload_data;
  wire ackNet_io_in_4_ready;
  wire ackNet_io_in_3_ready;
  wire ackNet_io_in_2_ready;
  wire ackNet_io_out_1_valid;
  wire[2:0] ackNet_io_out_1_bits_header_src;
  wire[2:0] ackNet_io_out_1_bits_header_dst;
  wire[3:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire ackNet_io_out_0_valid;
  wire[2:0] ackNet_io_out_0_bits_header_src;
  wire[2:0] ackNet_io_out_0_bits_header_dst;
  wire[3:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_io_client_release_ready;
  wire ClientTileLinkNetworkPort_io_network_acquire_valid;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_io_network_finish_valid;
  wire[2:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_io_network_release_valid;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_2_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_2_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_2_io_client_release_ready;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_valid;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_2_io_network_finish_valid;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire[3:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_2_io_network_release_valid;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire[5:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data;


  assign T0 = TileLinkEnqueuer_3_io_client_finish_ready;
  assign T1 = TileLinkEnqueuer_4_io_client_finish_ready;
  assign T2 = TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  assign T3 = TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  assign T4 = T5;
  assign T5 = TileLinkEnqueuer_io_manager_finish_bits_header_src + 3'h2;
  assign T6 = TileLinkEnqueuer_io_manager_finish_valid;
  assign T7 = TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  assign T8 = TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  assign T9 = T10;
  assign T10 = TileLinkEnqueuer_1_io_manager_finish_bits_header_src + 3'h2;
  assign T11 = TileLinkEnqueuer_1_io_manager_finish_valid;
  assign T12 = TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id;
  assign T13 = TileLinkEnqueuer_2_io_manager_finish_bits_header_dst;
  assign T14 = T15;
  assign T15 = TileLinkEnqueuer_2_io_manager_finish_bits_header_src + 3'h2;
  assign T16 = TileLinkEnqueuer_2_io_manager_finish_valid;
  assign T17 = TileLinkEnqueuer_io_manager_grant_ready;
  assign T18 = TileLinkEnqueuer_1_io_manager_grant_ready;
  assign T19 = TileLinkEnqueuer_2_io_manager_grant_ready;
  assign T20 = TileLinkEnqueuer_3_io_client_grant_bits_payload_data;
  assign T21 = TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type;
  assign T22 = TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type;
  assign T23 = TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id;
  assign T24 = TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id;
  assign T25 = TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat;
  assign T26 = T27;
  assign T27 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst + 3'h2;
  assign T28 = TileLinkEnqueuer_3_io_client_grant_bits_header_src;
  assign T29 = TileLinkEnqueuer_3_io_client_grant_valid;
  assign T30 = TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  assign T31 = TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  assign T32 = TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  assign T33 = TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  assign T34 = TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  assign T35 = TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  assign T36 = T37;
  assign T37 = TileLinkEnqueuer_4_io_client_grant_bits_header_dst + 3'h2;
  assign T38 = TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  assign T39 = TileLinkEnqueuer_4_io_client_grant_valid;
  assign T40 = TileLinkEnqueuer_io_manager_probe_ready;
  assign T41 = TileLinkEnqueuer_1_io_manager_probe_ready;
  assign T42 = TileLinkEnqueuer_2_io_manager_probe_ready;
  assign T43 = TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type;
  assign T44 = TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block;
  assign T45 = T46;
  assign T46 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst + 3'h2;
  assign T47 = TileLinkEnqueuer_3_io_client_probe_bits_header_src;
  assign T48 = TileLinkEnqueuer_3_io_client_probe_valid;
  assign T49 = TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  assign T50 = TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  assign T51 = T52;
  assign T52 = TileLinkEnqueuer_4_io_client_probe_bits_header_dst + 3'h2;
  assign T53 = TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  assign T54 = TileLinkEnqueuer_4_io_client_probe_valid;
  assign T55 = TileLinkEnqueuer_3_io_client_release_ready;
  assign T56 = TileLinkEnqueuer_4_io_client_release_ready;
  assign T57 = TileLinkEnqueuer_io_manager_release_bits_payload_data;
  assign T58 = TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  assign T59 = TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  assign T60 = TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  assign T61 = TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  assign T62 = TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  assign T63 = TileLinkEnqueuer_io_manager_release_bits_header_dst;
  assign T64 = T65;
  assign T65 = TileLinkEnqueuer_io_manager_release_bits_header_src + 3'h2;
  assign T66 = TileLinkEnqueuer_io_manager_release_valid;
  assign T67 = TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  assign T68 = TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  assign T69 = TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  assign T70 = TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  assign T71 = TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  assign T72 = TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  assign T73 = TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  assign T74 = T75;
  assign T75 = TileLinkEnqueuer_1_io_manager_release_bits_header_src + 3'h2;
  assign T76 = TileLinkEnqueuer_1_io_manager_release_valid;
  assign T77 = TileLinkEnqueuer_2_io_manager_release_bits_payload_data;
  assign T78 = TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type;
  assign T79 = TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary;
  assign T80 = TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id;
  assign T81 = TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block;
  assign T82 = TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat;
  assign T83 = TileLinkEnqueuer_2_io_manager_release_bits_header_dst;
  assign T84 = T85;
  assign T85 = TileLinkEnqueuer_2_io_manager_release_bits_header_src + 3'h2;
  assign T86 = TileLinkEnqueuer_2_io_manager_release_valid;
  assign T87 = TileLinkEnqueuer_3_io_client_acquire_ready;
  assign T88 = TileLinkEnqueuer_4_io_client_acquire_ready;
  assign T89 = TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  assign T90 = TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  assign T91 = TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  assign T92 = TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  assign T93 = TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  assign T94 = TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  assign T95 = TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  assign T96 = TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  assign T97 = T98;
  assign T98 = TileLinkEnqueuer_io_manager_acquire_bits_header_src + 3'h2;
  assign T99 = TileLinkEnqueuer_io_manager_acquire_valid;
  assign T100 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  assign T101 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  assign T102 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  assign T103 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign T104 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  assign T105 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  assign T106 = TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  assign T107 = TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  assign T108 = T109;
  assign T109 = TileLinkEnqueuer_1_io_manager_acquire_bits_header_src + 3'h2;
  assign T110 = TileLinkEnqueuer_1_io_manager_acquire_valid;
  assign T111 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data;
  assign T112 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union;
  assign T113 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type;
  assign T114 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type;
  assign T115 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat;
  assign T116 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id;
  assign T117 = TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block;
  assign T118 = TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst;
  assign T119 = T120;
  assign T120 = TileLinkEnqueuer_2_io_manager_acquire_bits_header_src + 3'h2;
  assign T121 = TileLinkEnqueuer_2_io_manager_acquire_valid;
  assign T122 = relNet_io_out_1_bits_payload_data;
  assign T123 = relNet_io_out_1_bits_payload_r_type;
  assign T124 = relNet_io_out_1_bits_payload_voluntary;
  assign T125 = relNet_io_out_1_bits_payload_client_xact_id;
  assign T126 = relNet_io_out_1_bits_payload_addr_block;
  assign T127 = relNet_io_out_1_bits_payload_addr_beat;
  assign T128 = relNet_io_out_1_bits_header_dst;
  assign T129 = T130;
  assign T130 = relNet_io_out_1_bits_header_src - 3'h2;
  assign T131 = relNet_io_out_1_valid;
  assign T132 = prbNet_io_in_1_ready;
  assign T133 = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T134 = ackNet_io_out_1_bits_header_dst;
  assign T135 = T136;
  assign T136 = ackNet_io_out_1_bits_header_src - 3'h2;
  assign T137 = ackNet_io_out_1_valid;
  assign T138 = gntNet_io_in_1_ready;
  assign T139 = acqNet_io_out_1_bits_payload_data;
  assign T140 = acqNet_io_out_1_bits_payload_union;
  assign T141 = acqNet_io_out_1_bits_payload_a_type;
  assign T142 = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T143 = acqNet_io_out_1_bits_payload_addr_beat;
  assign T144 = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T145 = acqNet_io_out_1_bits_payload_addr_block;
  assign T146 = acqNet_io_out_1_bits_header_dst;
  assign T147 = T148;
  assign T148 = acqNet_io_out_1_bits_header_src - 3'h2;
  assign T149 = acqNet_io_out_1_valid;
  assign T150 = relNet_io_out_0_bits_payload_data;
  assign T151 = relNet_io_out_0_bits_payload_r_type;
  assign T152 = relNet_io_out_0_bits_payload_voluntary;
  assign T153 = relNet_io_out_0_bits_payload_client_xact_id;
  assign T154 = relNet_io_out_0_bits_payload_addr_block;
  assign T155 = relNet_io_out_0_bits_payload_addr_beat;
  assign T156 = relNet_io_out_0_bits_header_dst;
  assign T157 = T158;
  assign T158 = relNet_io_out_0_bits_header_src - 3'h2;
  assign T159 = relNet_io_out_0_valid;
  assign T160 = prbNet_io_in_0_ready;
  assign T161 = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T162 = ackNet_io_out_0_bits_header_dst;
  assign T163 = T164;
  assign T164 = ackNet_io_out_0_bits_header_src - 3'h2;
  assign T165 = ackNet_io_out_0_valid;
  assign T166 = gntNet_io_in_0_ready;
  assign T167 = acqNet_io_out_0_bits_payload_data;
  assign T168 = acqNet_io_out_0_bits_payload_union;
  assign T169 = acqNet_io_out_0_bits_payload_a_type;
  assign T170 = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T171 = acqNet_io_out_0_bits_payload_addr_beat;
  assign T172 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T173 = acqNet_io_out_0_bits_payload_addr_block;
  assign T174 = acqNet_io_out_0_bits_header_dst;
  assign T175 = T176;
  assign T176 = acqNet_io_out_0_bits_header_src - 3'h2;
  assign T177 = acqNet_io_out_0_valid;
  assign T178 = relNet_io_in_4_ready;
  assign T179 = prbNet_io_out_4_bits_payload_p_type;
  assign T180 = prbNet_io_out_4_bits_payload_addr_block;
  assign T181 = T182;
  assign T182 = prbNet_io_out_4_bits_header_dst - 3'h2;
  assign T183 = prbNet_io_out_4_bits_header_src;
  assign T184 = prbNet_io_out_4_valid;
  assign T185 = ackNet_io_in_4_ready;
  assign T186 = gntNet_io_out_4_bits_payload_data;
  assign T187 = gntNet_io_out_4_bits_payload_g_type;
  assign T188 = gntNet_io_out_4_bits_payload_is_builtin_type;
  assign T189 = gntNet_io_out_4_bits_payload_manager_xact_id;
  assign T190 = gntNet_io_out_4_bits_payload_client_xact_id;
  assign T191 = gntNet_io_out_4_bits_payload_addr_beat;
  assign T192 = T193;
  assign T193 = gntNet_io_out_4_bits_header_dst - 3'h2;
  assign T194 = gntNet_io_out_4_bits_header_src;
  assign T195 = gntNet_io_out_4_valid;
  assign T196 = acqNet_io_in_4_ready;
  assign T197 = relNet_io_in_3_ready;
  assign T198 = prbNet_io_out_3_bits_payload_p_type;
  assign T199 = prbNet_io_out_3_bits_payload_addr_block;
  assign T200 = T201;
  assign T201 = prbNet_io_out_3_bits_header_dst - 3'h2;
  assign T202 = prbNet_io_out_3_bits_header_src;
  assign T203 = prbNet_io_out_3_valid;
  assign T204 = ackNet_io_in_3_ready;
  assign T205 = gntNet_io_out_3_bits_payload_data;
  assign T206 = gntNet_io_out_3_bits_payload_g_type;
  assign T207 = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T208 = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T209 = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T210 = gntNet_io_out_3_bits_payload_addr_beat;
  assign T211 = T212;
  assign T212 = gntNet_io_out_3_bits_header_dst - 3'h2;
  assign T213 = gntNet_io_out_3_bits_header_src;
  assign T214 = gntNet_io_out_3_valid;
  assign T215 = acqNet_io_in_3_ready;
  assign T216 = relNet_io_in_2_ready;
  assign T217 = prbNet_io_out_2_bits_payload_p_type;
  assign T218 = prbNet_io_out_2_bits_payload_addr_block;
  assign T219 = T220;
  assign T220 = prbNet_io_out_2_bits_header_dst - 3'h2;
  assign T221 = prbNet_io_out_2_bits_header_src;
  assign T222 = prbNet_io_out_2_valid;
  assign T223 = ackNet_io_in_2_ready;
  assign T224 = gntNet_io_out_2_bits_payload_data;
  assign T225 = gntNet_io_out_2_bits_payload_g_type;
  assign T226 = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T227 = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T228 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T229 = gntNet_io_out_2_bits_payload_addr_beat;
  assign T230 = T231;
  assign T231 = gntNet_io_out_2_bits_header_dst - 3'h2;
  assign T232 = gntNet_io_out_2_bits_header_src;
  assign T233 = gntNet_io_out_2_valid;
  assign T234 = acqNet_io_in_2_ready;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_io_manager_release_valid;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_io_manager_probe_ready;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_io_manager_finish_valid;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_io_manager_grant_ready;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_id;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_1_io_manager_release_bits_data;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_1_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_1_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_1_io_manager_release_valid;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_1_io_manager_probe_ready;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_1_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_1_io_manager_finish_valid;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_1_io_manager_grant_ready;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_id;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_1_io_manager_acquire_valid;
  assign io_clients_0_release_ready = ClientTileLinkNetworkPort_io_client_release_ready;
  assign io_clients_0_probe_bits_p_type = ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  assign io_clients_0_probe_bits_addr_block = ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  assign io_clients_0_probe_valid = ClientTileLinkNetworkPort_io_client_probe_valid;
  assign io_clients_0_grant_bits_data = ClientTileLinkNetworkPort_io_client_grant_bits_data;
  assign io_clients_0_grant_bits_g_type = ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  assign io_clients_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  assign io_clients_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  assign io_clients_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  assign io_clients_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  assign io_clients_0_grant_valid = ClientTileLinkNetworkPort_io_client_grant_valid;
  assign io_clients_0_acquire_ready = ClientTileLinkNetworkPort_io_client_acquire_ready;
  assign io_clients_1_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_1_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_1_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_1_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_1_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_1_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_1_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_1_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_1_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_1_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_1_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_1_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_2_release_ready = ClientTileLinkNetworkPort_2_io_client_release_ready;
  assign io_clients_2_probe_bits_p_type = ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  assign io_clients_2_probe_bits_addr_block = ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  assign io_clients_2_probe_valid = ClientTileLinkNetworkPort_2_io_client_probe_valid;
  assign io_clients_2_grant_bits_data = ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  assign io_clients_2_grant_bits_g_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  assign io_clients_2_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  assign io_clients_2_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  assign io_clients_2_grant_bits_client_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  assign io_clients_2_grant_bits_addr_beat = ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  assign io_clients_2_grant_valid = ClientTileLinkNetworkPort_2_io_client_grant_valid;
  assign io_clients_2_acquire_ready = ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  ClientTileLinkNetworkPort_0 ClientTileLinkNetworkPort(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_0_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_0_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_0_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_0_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_0_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_0_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_0_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_0_acquire_bits_data ),
       .io_client_grant_ready( io_clients_0_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_0_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_io_client_release_ready ),
       .io_client_release_valid( io_clients_0_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_0_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_0_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_0_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_0_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_0_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_0_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( T234 ),
       .io_manager_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_manager_grant_valid( T233 ),
       .io_manager_grant_bits_header_src( T232 ),
       .io_manager_grant_bits_header_dst( T230 ),
       .io_manager_grant_bits_payload_addr_beat( T229 ),
       .io_manager_grant_bits_payload_client_xact_id( T228 ),
       .io_manager_grant_bits_payload_manager_xact_id( T227 ),
       .io_manager_grant_bits_payload_is_builtin_type( T226 ),
       .io_manager_grant_bits_payload_g_type( T225 ),
       .io_manager_grant_bits_payload_data( T224 ),
       .io_manager_finish_ready( T223 ),
       .io_manager_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_manager_probe_valid( T222 ),
       .io_manager_probe_bits_header_src( T221 ),
       .io_manager_probe_bits_header_dst( T219 ),
       .io_manager_probe_bits_payload_addr_block( T218 ),
       .io_manager_probe_bits_payload_p_type( T217 ),
       .io_manager_release_ready( T216 ),
       .io_manager_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_1 ClientTileLinkNetworkPort_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_1_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_1_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_1_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_1_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_1_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_1_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_1_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_1_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_1_acquire_bits_data ),
       .io_client_grant_ready( io_clients_1_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_1_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_1_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_1_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_1_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_1_io_client_release_ready ),
       .io_client_release_valid( io_clients_1_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_1_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_1_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_1_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_1_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_1_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_1_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( T215 ),
       .io_manager_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_manager_grant_valid( T214 ),
       .io_manager_grant_bits_header_src( T213 ),
       .io_manager_grant_bits_header_dst( T211 ),
       .io_manager_grant_bits_payload_addr_beat( T210 ),
       .io_manager_grant_bits_payload_client_xact_id( T209 ),
       .io_manager_grant_bits_payload_manager_xact_id( T208 ),
       .io_manager_grant_bits_payload_is_builtin_type( T207 ),
       .io_manager_grant_bits_payload_g_type( T206 ),
       .io_manager_grant_bits_payload_data( T205 ),
       .io_manager_finish_ready( T204 ),
       .io_manager_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_manager_probe_valid( T203 ),
       .io_manager_probe_bits_header_src( T202 ),
       .io_manager_probe_bits_header_dst( T200 ),
       .io_manager_probe_bits_payload_addr_block( T199 ),
       .io_manager_probe_bits_payload_p_type( T198 ),
       .io_manager_release_ready( T197 ),
       .io_manager_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_2 ClientTileLinkNetworkPort_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_2_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_2_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_2_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_2_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_2_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_2_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_2_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_2_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_2_acquire_bits_data ),
       .io_client_grant_ready( io_clients_2_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_2_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_2_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_2_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_2_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_2_io_client_release_ready ),
       .io_client_release_valid( io_clients_2_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_2_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_2_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_2_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_2_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_2_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_2_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( T196 ),
       .io_manager_acquire_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_2_io_manager_grant_ready ),
       .io_manager_grant_valid( T195 ),
       .io_manager_grant_bits_header_src( T194 ),
       .io_manager_grant_bits_header_dst( T192 ),
       .io_manager_grant_bits_payload_addr_beat( T191 ),
       .io_manager_grant_bits_payload_client_xact_id( T190 ),
       .io_manager_grant_bits_payload_manager_xact_id( T189 ),
       .io_manager_grant_bits_payload_is_builtin_type( T188 ),
       .io_manager_grant_bits_payload_g_type( T187 ),
       .io_manager_grant_bits_payload_data( T186 ),
       .io_manager_finish_ready( T185 ),
       .io_manager_finish_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_2_io_manager_probe_ready ),
       .io_manager_probe_valid( T184 ),
       .io_manager_probe_bits_header_src( T183 ),
       .io_manager_probe_bits_header_dst( T181 ),
       .io_manager_probe_bits_payload_addr_block( T180 ),
       .io_manager_probe_bits_payload_p_type( T179 ),
       .io_manager_release_ready( T178 ),
       .io_manager_release_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data )
  );
  ManagerTileLinkNetworkPort_0 ManagerTileLinkNetworkPort(
       .io_manager_acquire_ready( io_managers_0_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_0_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_0_grant_bits_addr_beat ),
       .io_manager_grant_bits_client_xact_id( io_managers_0_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_0_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_0_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_0_grant_bits_g_type ),
       .io_manager_grant_bits_data( io_managers_0_grant_bits_data ),
       .io_manager_grant_bits_client_id( io_managers_0_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_0_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_0_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_0_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_0_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_0_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_0_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_io_manager_release_valid ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_io_manager_release_bits_r_type ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_io_manager_release_bits_data ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_network_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_3(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_client_acquire_valid( T177 ),
       .io_client_acquire_bits_header_src( T175 ),
       .io_client_acquire_bits_header_dst( T174 ),
       .io_client_acquire_bits_payload_addr_block( T173 ),
       .io_client_acquire_bits_payload_client_xact_id( T172 ),
       .io_client_acquire_bits_payload_addr_beat( T171 ),
       .io_client_acquire_bits_payload_is_builtin_type( T170 ),
       .io_client_acquire_bits_payload_a_type( T169 ),
       .io_client_acquire_bits_payload_union( T168 ),
       .io_client_acquire_bits_payload_data( T167 ),
       .io_client_grant_ready( T166 ),
       .io_client_grant_valid( TileLinkEnqueuer_3_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_client_finish_valid( T165 ),
       .io_client_finish_bits_header_src( T163 ),
       .io_client_finish_bits_header_dst( T162 ),
       .io_client_finish_bits_payload_manager_xact_id( T161 ),
       .io_client_probe_ready( T160 ),
       .io_client_probe_valid( TileLinkEnqueuer_3_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_client_release_valid( T159 ),
       .io_client_release_bits_header_src( T157 ),
       .io_client_release_bits_header_dst( T156 ),
       .io_client_release_bits_payload_addr_beat( T155 ),
       .io_client_release_bits_payload_addr_block( T154 ),
       .io_client_release_bits_payload_client_xact_id( T153 ),
       .io_client_release_bits_payload_voluntary( T152 ),
       .io_client_release_bits_payload_r_type( T151 ),
       .io_client_release_bits_payload_data( T150 ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort_1(
       .io_manager_acquire_ready( io_managers_1_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_1_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_1_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_1_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_1_grant_bits_addr_beat ),
       .io_manager_grant_bits_client_xact_id( io_managers_1_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_1_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_1_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_1_grant_bits_g_type ),
       .io_manager_grant_bits_data( io_managers_1_grant_bits_data ),
       .io_manager_grant_bits_client_id( io_managers_1_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_1_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_1_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_1_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_1_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_1_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_1_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_1_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_1_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_1_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_1_io_manager_release_valid ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_1_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_1_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_1_io_manager_release_bits_r_type ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_1_io_manager_release_bits_data ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_1_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_1_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_4_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_4_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data ),
       .io_network_grant_ready( TileLinkEnqueuer_4_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_1_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_data ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_1_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_4_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_4_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_4_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_4_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_1_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_1_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_4_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_4_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_4_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_4_io_manager_release_bits_payload_data )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_4(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_4_io_client_acquire_ready ),
       .io_client_acquire_valid( T149 ),
       .io_client_acquire_bits_header_src( T147 ),
       .io_client_acquire_bits_header_dst( T146 ),
       .io_client_acquire_bits_payload_addr_block( T145 ),
       .io_client_acquire_bits_payload_client_xact_id( T144 ),
       .io_client_acquire_bits_payload_addr_beat( T143 ),
       .io_client_acquire_bits_payload_is_builtin_type( T142 ),
       .io_client_acquire_bits_payload_a_type( T141 ),
       .io_client_acquire_bits_payload_union( T140 ),
       .io_client_acquire_bits_payload_data( T139 ),
       .io_client_grant_ready( T138 ),
       .io_client_grant_valid( TileLinkEnqueuer_4_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_4_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_4_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_4_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_4_io_client_finish_ready ),
       .io_client_finish_valid( T137 ),
       .io_client_finish_bits_header_src( T135 ),
       .io_client_finish_bits_header_dst( T134 ),
       .io_client_finish_bits_payload_manager_xact_id( T133 ),
       .io_client_probe_ready( T132 ),
       .io_client_probe_valid( TileLinkEnqueuer_4_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_4_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_4_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_4_io_client_release_ready ),
       .io_client_release_valid( T131 ),
       .io_client_release_bits_header_src( T129 ),
       .io_client_release_bits_header_dst( T128 ),
       .io_client_release_bits_payload_addr_beat( T127 ),
       .io_client_release_bits_payload_addr_block( T126 ),
       .io_client_release_bits_payload_client_xact_id( T125 ),
       .io_client_release_bits_payload_voluntary( T124 ),
       .io_client_release_bits_payload_r_type( T123 ),
       .io_client_release_bits_payload_data( T122 ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_1_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_4_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_4_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_4_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_1_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_1_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_1_io_network_grant_bits_payload_data ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_1_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_4_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_4_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_4_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_4_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_1_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_1_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_1_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_4_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_4_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_4_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_4_io_manager_release_bits_payload_data )
  );
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_4_ready( acqNet_io_in_4_ready ),
       .io_in_4_valid( T121 ),
       .io_in_4_bits_header_src( T119 ),
       .io_in_4_bits_header_dst( T118 ),
       .io_in_4_bits_payload_addr_block( T117 ),
       .io_in_4_bits_payload_client_xact_id( T116 ),
       .io_in_4_bits_payload_addr_beat( T115 ),
       .io_in_4_bits_payload_is_builtin_type( T114 ),
       .io_in_4_bits_payload_a_type( T113 ),
       .io_in_4_bits_payload_union( T112 ),
       .io_in_4_bits_payload_data( T111 ),
       .io_in_3_ready( acqNet_io_in_3_ready ),
       .io_in_3_valid( T110 ),
       .io_in_3_bits_header_src( T108 ),
       .io_in_3_bits_header_dst( T107 ),
       .io_in_3_bits_payload_addr_block( T106 ),
       .io_in_3_bits_payload_client_xact_id( T105 ),
       .io_in_3_bits_payload_addr_beat( T104 ),
       .io_in_3_bits_payload_is_builtin_type( T103 ),
       .io_in_3_bits_payload_a_type( T102 ),
       .io_in_3_bits_payload_union( T101 ),
       .io_in_3_bits_payload_data( T100 ),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T99 ),
       .io_in_2_bits_header_src( T97 ),
       .io_in_2_bits_header_dst( T96 ),
       .io_in_2_bits_payload_addr_block( T95 ),
       .io_in_2_bits_payload_client_xact_id( T94 ),
       .io_in_2_bits_payload_addr_beat( T93 ),
       .io_in_2_bits_payload_is_builtin_type( T92 ),
       .io_in_2_bits_payload_a_type( T91 ),
       .io_in_2_bits_payload_union( T90 ),
       .io_in_2_bits_payload_data( T89 ),
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr_block(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_addr_beat(  )
       //.io_in_1_bits_payload_is_builtin_type(  )
       //.io_in_1_bits_payload_a_type(  )
       //.io_in_1_bits_payload_union(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr_block(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_addr_beat(  )
       //.io_in_0_bits_payload_is_builtin_type(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_union(  )
       //.io_in_0_bits_payload_data(  )
       .io_out_4_ready( 1'h0 ),
       //.io_out_4_valid(  )
       //.io_out_4_bits_header_src(  )
       //.io_out_4_bits_header_dst(  )
       //.io_out_4_bits_payload_addr_block(  )
       //.io_out_4_bits_payload_client_xact_id(  )
       //.io_out_4_bits_payload_addr_beat(  )
       //.io_out_4_bits_payload_is_builtin_type(  )
       //.io_out_4_bits_payload_a_type(  )
       //.io_out_4_bits_payload_union(  )
       //.io_out_4_bits_payload_data(  )
       .io_out_3_ready( 1'h0 ),
       //.io_out_3_valid(  )
       //.io_out_3_bits_header_src(  )
       //.io_out_3_bits_header_dst(  )
       //.io_out_3_bits_payload_addr_block(  )
       //.io_out_3_bits_payload_client_xact_id(  )
       //.io_out_3_bits_payload_addr_beat(  )
       //.io_out_3_bits_payload_is_builtin_type(  )
       //.io_out_3_bits_payload_a_type(  )
       //.io_out_3_bits_payload_union(  )
       //.io_out_3_bits_payload_data(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr_block(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_addr_beat(  )
       //.io_out_2_bits_payload_is_builtin_type(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_union(  )
       //.io_out_2_bits_payload_data(  )
       .io_out_1_ready( T88 ),
       .io_out_1_valid( acqNet_io_out_1_valid ),
       .io_out_1_bits_header_src( acqNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( acqNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr_block( acqNet_io_out_1_bits_payload_addr_block ),
       .io_out_1_bits_payload_client_xact_id( acqNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_addr_beat( acqNet_io_out_1_bits_payload_addr_beat ),
       .io_out_1_bits_payload_is_builtin_type( acqNet_io_out_1_bits_payload_is_builtin_type ),
       .io_out_1_bits_payload_a_type( acqNet_io_out_1_bits_payload_a_type ),
       .io_out_1_bits_payload_union( acqNet_io_out_1_bits_payload_union ),
       .io_out_1_bits_payload_data( acqNet_io_out_1_bits_payload_data ),
       .io_out_0_ready( T87 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr_block( acqNet_io_out_0_bits_payload_addr_block ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_addr_beat( acqNet_io_out_0_bits_payload_addr_beat ),
       .io_out_0_bits_payload_is_builtin_type( acqNet_io_out_0_bits_payload_is_builtin_type ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_union( acqNet_io_out_0_bits_payload_union ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign acqNet.io_in_1_bits_header_src = {1{$random}};
    assign acqNet.io_in_1_bits_header_dst = {1{$random}};
    assign acqNet.io_in_1_bits_payload_addr_block = {1{$random}};
    assign acqNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_1_bits_payload_addr_beat = {1{$random}};
    assign acqNet.io_in_1_bits_payload_is_builtin_type = {1{$random}};
    assign acqNet.io_in_1_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_1_bits_payload_union = {1{$random}};
    assign acqNet.io_in_1_bits_payload_data = {4{$random}};
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr_block = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr_beat = {1{$random}};
    assign acqNet.io_in_0_bits_payload_is_builtin_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_union = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {4{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_4_ready( relNet_io_in_4_ready ),
       .io_in_4_valid( T86 ),
       .io_in_4_bits_header_src( T84 ),
       .io_in_4_bits_header_dst( T83 ),
       .io_in_4_bits_payload_addr_beat( T82 ),
       .io_in_4_bits_payload_addr_block( T81 ),
       .io_in_4_bits_payload_client_xact_id( T80 ),
       .io_in_4_bits_payload_voluntary( T79 ),
       .io_in_4_bits_payload_r_type( T78 ),
       .io_in_4_bits_payload_data( T77 ),
       .io_in_3_ready( relNet_io_in_3_ready ),
       .io_in_3_valid( T76 ),
       .io_in_3_bits_header_src( T74 ),
       .io_in_3_bits_header_dst( T73 ),
       .io_in_3_bits_payload_addr_beat( T72 ),
       .io_in_3_bits_payload_addr_block( T71 ),
       .io_in_3_bits_payload_client_xact_id( T70 ),
       .io_in_3_bits_payload_voluntary( T69 ),
       .io_in_3_bits_payload_r_type( T68 ),
       .io_in_3_bits_payload_data( T67 ),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T66 ),
       .io_in_2_bits_header_src( T64 ),
       .io_in_2_bits_header_dst( T63 ),
       .io_in_2_bits_payload_addr_beat( T62 ),
       .io_in_2_bits_payload_addr_block( T61 ),
       .io_in_2_bits_payload_client_xact_id( T60 ),
       .io_in_2_bits_payload_voluntary( T59 ),
       .io_in_2_bits_payload_r_type( T58 ),
       .io_in_2_bits_payload_data( T57 ),
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr_beat(  )
       //.io_in_1_bits_payload_addr_block(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_voluntary(  )
       //.io_in_1_bits_payload_r_type(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr_beat(  )
       //.io_in_0_bits_payload_addr_block(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_voluntary(  )
       //.io_in_0_bits_payload_r_type(  )
       //.io_in_0_bits_payload_data(  )
       .io_out_4_ready( 1'h0 ),
       //.io_out_4_valid(  )
       //.io_out_4_bits_header_src(  )
       //.io_out_4_bits_header_dst(  )
       //.io_out_4_bits_payload_addr_beat(  )
       //.io_out_4_bits_payload_addr_block(  )
       //.io_out_4_bits_payload_client_xact_id(  )
       //.io_out_4_bits_payload_voluntary(  )
       //.io_out_4_bits_payload_r_type(  )
       //.io_out_4_bits_payload_data(  )
       .io_out_3_ready( 1'h0 ),
       //.io_out_3_valid(  )
       //.io_out_3_bits_header_src(  )
       //.io_out_3_bits_header_dst(  )
       //.io_out_3_bits_payload_addr_beat(  )
       //.io_out_3_bits_payload_addr_block(  )
       //.io_out_3_bits_payload_client_xact_id(  )
       //.io_out_3_bits_payload_voluntary(  )
       //.io_out_3_bits_payload_r_type(  )
       //.io_out_3_bits_payload_data(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr_beat(  )
       //.io_out_2_bits_payload_addr_block(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_voluntary(  )
       //.io_out_2_bits_payload_r_type(  )
       //.io_out_2_bits_payload_data(  )
       .io_out_1_ready( T56 ),
       .io_out_1_valid( relNet_io_out_1_valid ),
       .io_out_1_bits_header_src( relNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( relNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr_beat( relNet_io_out_1_bits_payload_addr_beat ),
       .io_out_1_bits_payload_addr_block( relNet_io_out_1_bits_payload_addr_block ),
       .io_out_1_bits_payload_client_xact_id( relNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_voluntary( relNet_io_out_1_bits_payload_voluntary ),
       .io_out_1_bits_payload_r_type( relNet_io_out_1_bits_payload_r_type ),
       .io_out_1_bits_payload_data( relNet_io_out_1_bits_payload_data ),
       .io_out_0_ready( T55 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr_beat( relNet_io_out_0_bits_payload_addr_beat ),
       .io_out_0_bits_payload_addr_block( relNet_io_out_0_bits_payload_addr_block ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_voluntary( relNet_io_out_0_bits_payload_voluntary ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign relNet.io_in_1_bits_header_src = {1{$random}};
    assign relNet.io_in_1_bits_header_dst = {1{$random}};
    assign relNet.io_in_1_bits_payload_addr_beat = {1{$random}};
    assign relNet.io_in_1_bits_payload_addr_block = {1{$random}};
    assign relNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_1_bits_payload_voluntary = {1{$random}};
    assign relNet.io_in_1_bits_payload_r_type = {1{$random}};
    assign relNet.io_in_1_bits_payload_data = {4{$random}};
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr_beat = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr_block = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_voluntary = {1{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {4{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_4_ready(  )
       .io_in_4_valid( 1'h0 ),
       //.io_in_4_bits_header_src(  )
       //.io_in_4_bits_header_dst(  )
       //.io_in_4_bits_payload_addr_block(  )
       //.io_in_4_bits_payload_p_type(  )
       //.io_in_3_ready(  )
       .io_in_3_valid( 1'h0 ),
       //.io_in_3_bits_header_src(  )
       //.io_in_3_bits_header_dst(  )
       //.io_in_3_bits_payload_addr_block(  )
       //.io_in_3_bits_payload_p_type(  )
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr_block(  )
       //.io_in_2_bits_payload_p_type(  )
       .io_in_1_ready( prbNet_io_in_1_ready ),
       .io_in_1_valid( T54 ),
       .io_in_1_bits_header_src( T53 ),
       .io_in_1_bits_header_dst( T51 ),
       .io_in_1_bits_payload_addr_block( T50 ),
       .io_in_1_bits_payload_p_type( T49 ),
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T48 ),
       .io_in_0_bits_header_src( T47 ),
       .io_in_0_bits_header_dst( T45 ),
       .io_in_0_bits_payload_addr_block( T44 ),
       .io_in_0_bits_payload_p_type( T43 ),
       .io_out_4_ready( T42 ),
       .io_out_4_valid( prbNet_io_out_4_valid ),
       .io_out_4_bits_header_src( prbNet_io_out_4_bits_header_src ),
       .io_out_4_bits_header_dst( prbNet_io_out_4_bits_header_dst ),
       .io_out_4_bits_payload_addr_block( prbNet_io_out_4_bits_payload_addr_block ),
       .io_out_4_bits_payload_p_type( prbNet_io_out_4_bits_payload_p_type ),
       .io_out_3_ready( T41 ),
       .io_out_3_valid( prbNet_io_out_3_valid ),
       .io_out_3_bits_header_src( prbNet_io_out_3_bits_header_src ),
       .io_out_3_bits_header_dst( prbNet_io_out_3_bits_header_dst ),
       .io_out_3_bits_payload_addr_block( prbNet_io_out_3_bits_payload_addr_block ),
       .io_out_3_bits_payload_p_type( prbNet_io_out_3_bits_payload_p_type ),
       .io_out_2_ready( T40 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr_block( prbNet_io_out_2_bits_payload_addr_block ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr_block(  )
       //.io_out_1_bits_payload_p_type(  )
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr_block(  )
       //.io_out_0_bits_payload_p_type(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign prbNet.io_in_4_bits_header_src = {1{$random}};
    assign prbNet.io_in_4_bits_header_dst = {1{$random}};
    assign prbNet.io_in_4_bits_payload_addr_block = {1{$random}};
    assign prbNet.io_in_4_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_3_bits_header_src = {1{$random}};
    assign prbNet.io_in_3_bits_header_dst = {1{$random}};
    assign prbNet.io_in_3_bits_payload_addr_block = {1{$random}};
    assign prbNet.io_in_3_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr_block = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_4_ready(  )
       .io_in_4_valid( 1'h0 ),
       //.io_in_4_bits_header_src(  )
       //.io_in_4_bits_header_dst(  )
       //.io_in_4_bits_payload_addr_beat(  )
       //.io_in_4_bits_payload_client_xact_id(  )
       //.io_in_4_bits_payload_manager_xact_id(  )
       //.io_in_4_bits_payload_is_builtin_type(  )
       //.io_in_4_bits_payload_g_type(  )
       //.io_in_4_bits_payload_data(  )
       //.io_in_3_ready(  )
       .io_in_3_valid( 1'h0 ),
       //.io_in_3_bits_header_src(  )
       //.io_in_3_bits_header_dst(  )
       //.io_in_3_bits_payload_addr_beat(  )
       //.io_in_3_bits_payload_client_xact_id(  )
       //.io_in_3_bits_payload_manager_xact_id(  )
       //.io_in_3_bits_payload_is_builtin_type(  )
       //.io_in_3_bits_payload_g_type(  )
       //.io_in_3_bits_payload_data(  )
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr_beat(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_manager_xact_id(  )
       //.io_in_2_bits_payload_is_builtin_type(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_2_bits_payload_data(  )
       .io_in_1_ready( gntNet_io_in_1_ready ),
       .io_in_1_valid( T39 ),
       .io_in_1_bits_header_src( T38 ),
       .io_in_1_bits_header_dst( T36 ),
       .io_in_1_bits_payload_addr_beat( T35 ),
       .io_in_1_bits_payload_client_xact_id( T34 ),
       .io_in_1_bits_payload_manager_xact_id( T33 ),
       .io_in_1_bits_payload_is_builtin_type( T32 ),
       .io_in_1_bits_payload_g_type( T31 ),
       .io_in_1_bits_payload_data( T30 ),
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T29 ),
       .io_in_0_bits_header_src( T28 ),
       .io_in_0_bits_header_dst( T26 ),
       .io_in_0_bits_payload_addr_beat( T25 ),
       .io_in_0_bits_payload_client_xact_id( T24 ),
       .io_in_0_bits_payload_manager_xact_id( T23 ),
       .io_in_0_bits_payload_is_builtin_type( T22 ),
       .io_in_0_bits_payload_g_type( T21 ),
       .io_in_0_bits_payload_data( T20 ),
       .io_out_4_ready( T19 ),
       .io_out_4_valid( gntNet_io_out_4_valid ),
       .io_out_4_bits_header_src( gntNet_io_out_4_bits_header_src ),
       .io_out_4_bits_header_dst( gntNet_io_out_4_bits_header_dst ),
       .io_out_4_bits_payload_addr_beat( gntNet_io_out_4_bits_payload_addr_beat ),
       .io_out_4_bits_payload_client_xact_id( gntNet_io_out_4_bits_payload_client_xact_id ),
       .io_out_4_bits_payload_manager_xact_id( gntNet_io_out_4_bits_payload_manager_xact_id ),
       .io_out_4_bits_payload_is_builtin_type( gntNet_io_out_4_bits_payload_is_builtin_type ),
       .io_out_4_bits_payload_g_type( gntNet_io_out_4_bits_payload_g_type ),
       .io_out_4_bits_payload_data( gntNet_io_out_4_bits_payload_data ),
       .io_out_3_ready( T18 ),
       .io_out_3_valid( gntNet_io_out_3_valid ),
       .io_out_3_bits_header_src( gntNet_io_out_3_bits_header_src ),
       .io_out_3_bits_header_dst( gntNet_io_out_3_bits_header_dst ),
       .io_out_3_bits_payload_addr_beat( gntNet_io_out_3_bits_payload_addr_beat ),
       .io_out_3_bits_payload_client_xact_id( gntNet_io_out_3_bits_payload_client_xact_id ),
       .io_out_3_bits_payload_manager_xact_id( gntNet_io_out_3_bits_payload_manager_xact_id ),
       .io_out_3_bits_payload_is_builtin_type( gntNet_io_out_3_bits_payload_is_builtin_type ),
       .io_out_3_bits_payload_g_type( gntNet_io_out_3_bits_payload_g_type ),
       .io_out_3_bits_payload_data( gntNet_io_out_3_bits_payload_data ),
       .io_out_2_ready( T17 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr_beat( gntNet_io_out_2_bits_payload_addr_beat ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_manager_xact_id( gntNet_io_out_2_bits_payload_manager_xact_id ),
       .io_out_2_bits_payload_is_builtin_type( gntNet_io_out_2_bits_payload_is_builtin_type ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr_beat(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_manager_xact_id(  )
       //.io_out_1_bits_payload_is_builtin_type(  )
       //.io_out_1_bits_payload_g_type(  )
       //.io_out_1_bits_payload_data(  )
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr_beat(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_manager_xact_id(  )
       //.io_out_0_bits_payload_is_builtin_type(  )
       //.io_out_0_bits_payload_g_type(  )
       //.io_out_0_bits_payload_data(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign gntNet.io_in_4_bits_header_src = {1{$random}};
    assign gntNet.io_in_4_bits_header_dst = {1{$random}};
    assign gntNet.io_in_4_bits_payload_addr_beat = {1{$random}};
    assign gntNet.io_in_4_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_4_bits_payload_manager_xact_id = {1{$random}};
    assign gntNet.io_in_4_bits_payload_is_builtin_type = {1{$random}};
    assign gntNet.io_in_4_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_4_bits_payload_data = {4{$random}};
    assign gntNet.io_in_3_bits_header_src = {1{$random}};
    assign gntNet.io_in_3_bits_header_dst = {1{$random}};
    assign gntNet.io_in_3_bits_payload_addr_beat = {1{$random}};
    assign gntNet.io_in_3_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_3_bits_payload_manager_xact_id = {1{$random}};
    assign gntNet.io_in_3_bits_payload_is_builtin_type = {1{$random}};
    assign gntNet.io_in_3_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_3_bits_payload_data = {4{$random}};
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_addr_beat = {1{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_manager_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_is_builtin_type = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {4{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_4_ready( ackNet_io_in_4_ready ),
       .io_in_4_valid( T16 ),
       .io_in_4_bits_header_src( T14 ),
       .io_in_4_bits_header_dst( T13 ),
       .io_in_4_bits_payload_manager_xact_id( T12 ),
       .io_in_3_ready( ackNet_io_in_3_ready ),
       .io_in_3_valid( T11 ),
       .io_in_3_bits_header_src( T9 ),
       .io_in_3_bits_header_dst( T8 ),
       .io_in_3_bits_payload_manager_xact_id( T7 ),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T6 ),
       .io_in_2_bits_header_src( T4 ),
       .io_in_2_bits_header_dst( T3 ),
       .io_in_2_bits_payload_manager_xact_id( T2 ),
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_manager_xact_id(  )
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_manager_xact_id(  )
       .io_out_4_ready( 1'h0 ),
       //.io_out_4_valid(  )
       //.io_out_4_bits_header_src(  )
       //.io_out_4_bits_header_dst(  )
       //.io_out_4_bits_payload_manager_xact_id(  )
       .io_out_3_ready( 1'h0 ),
       //.io_out_3_valid(  )
       //.io_out_3_bits_header_src(  )
       //.io_out_3_bits_header_dst(  )
       //.io_out_3_bits_payload_manager_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_manager_xact_id(  )
       .io_out_1_ready( T1 ),
       .io_out_1_valid( ackNet_io_out_1_valid ),
       .io_out_1_bits_header_src( ackNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( ackNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_manager_xact_id( ackNet_io_out_1_bits_payload_manager_xact_id ),
       .io_out_0_ready( T0 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_manager_xact_id( ackNet_io_out_0_bits_payload_manager_xact_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ackNet.io_in_1_bits_header_src = {1{$random}};
    assign ackNet.io_in_1_bits_header_dst = {1{$random}};
    assign ackNet.io_in_1_bits_payload_manager_xact_id = {1{$random}};
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_manager_xact_id = {1{$random}};
// synthesis translate_on
`endif
endmodule

module BroadcastVoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[25:0] io_inner_probe_bits_addr_block
    //output[1:0] io_inner_probe_bits_p_type
    //output[1:0] io_inner_probe_bits_client_id
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  state;
  wire T148;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire all_pending_done;
  wire T14;
  reg  pending_ignt;
  wire T149;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [3:0] pending_writes;
  wire[3:0] T150;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T151;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[3:0] T36;
  wire[3:0] T37;
  wire[3:0] T152;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[3:0] T48;
  wire[3:0] T153;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  reg [3:0] pending_irels;
  wire[3:0] T154;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T155;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[3:0] T74;
  wire[3:0] T75;
  wire[3:0] T76;
  wire[3:0] T156;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] T97;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire[1:0] T102;
  wire T103;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[1:0] T108;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire T160;
  wire T161;
  wire T162;
  wire[3:0] T109;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T110;
  wire T111;
  wire T112;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[16:0] T118;
  wire[16:0] T119;
  wire[15:0] T120;
  wire[2:0] T121;
  wire T122;
  wire[1:0] T123;
  wire[3:0] T163;
  wire[5:0] T124;
  wire[25:0] T125;
  reg [25:0] xact_addr_block;
  wire[25:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[1:0] T134;
  reg [1:0] xact_client_id;
  wire[1:0] T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire T138;
  wire[3:0] T139;
  wire[5:0] T140;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    pending_ignt = {1{$random}};
    pending_writes = {1{$random}};
    pending_irels = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_addr_block = {1{$random}};
    xact_client_id = {1{$random}};
    xact_client_xact_id = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_inner_probe_bits_client_id = {1{$random}};
//  assign io_inner_probe_bits_p_type = {1{$random}};
//  assign io_inner_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T5 = T7 & T6;
  assign T6 = io_inner_release_ready & io_inner_release_valid;
  assign T7 = state == 1'h0;
  assign T148 = reset ? 1'h0 : T8;
  assign T8 = T13 ? 1'h0 : T9;
  assign T9 = T10 ? 1'h1 : state;
  assign T10 = T12 & T11;
  assign T11 = io_inner_release_ready & io_inner_release_valid;
  assign T12 = state == 1'h0;
  assign T13 = T92 & all_pending_done;
  assign all_pending_done = T14 ^ 1'h1;
  assign T14 = T18 | pending_ignt;
  assign T149 = reset ? 1'h0 : T15;
  assign T15 = T10 ? 1'h1 : T16;
  assign T16 = T17 ? 1'h0 : pending_ignt;
  assign T17 = io_inner_grant_ready & io_inner_grant_valid;
  assign T18 = T56 | T19;
  assign T19 = pending_writes != 4'h0;
  assign T150 = reset ? 4'h0 : T20;
  assign T20 = T10 ? T46 : T21;
  assign T21 = T32 | T22;
  assign T22 = T24 & T23;
  assign T23 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T24 = 4'h0 - T151;
  assign T151 = {3'h0, T25};
  assign T25 = T31 & T26;
  assign T26 = T28 | T27;
  assign T27 = 3'h2 == io_inner_release_bits_r_type;
  assign T28 = T30 | T29;
  assign T29 = 3'h1 == io_inner_release_bits_r_type;
  assign T30 = 3'h0 == io_inner_release_bits_r_type;
  assign T31 = io_inner_release_ready & io_inner_release_valid;
  assign T32 = pending_writes & T33;
  assign T33 = T36 | T34;
  assign T34 = ~ T35;
  assign T35 = 1'h1 << io_outer_acquire_bits_addr_beat;
  assign T36 = ~ T37;
  assign T37 = 4'h0 - T152;
  assign T152 = {3'h0, T38};
  assign T38 = T45 & T39;
  assign T39 = io_outer_acquire_bits_is_builtin_type & T40;
  assign T40 = T42 | T41;
  assign T41 = 3'h4 == io_outer_acquire_bits_a_type;
  assign T42 = T44 | T43;
  assign T43 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T44 = 3'h2 == io_outer_acquire_bits_a_type;
  assign T45 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T46 = T48 & T47;
  assign T47 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T48 = 4'h0 - T153;
  assign T153 = {3'h0, T49};
  assign T49 = T55 & T50;
  assign T50 = T52 | T51;
  assign T51 = 3'h2 == io_inner_release_bits_r_type;
  assign T52 = T54 | T53;
  assign T53 = 3'h1 == io_inner_release_bits_r_type;
  assign T54 = 3'h0 == io_inner_release_bits_r_type;
  assign T55 = io_inner_release_ready & io_inner_release_valid;
  assign T56 = pending_irels != 4'h0;
  assign T154 = reset ? 4'h0 : T57;
  assign T57 = T90 ? 4'h0 : T58;
  assign T58 = T84 ? T72 : T59;
  assign T59 = pending_irels & T60;
  assign T60 = T63 | T61;
  assign T61 = ~ T62;
  assign T62 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T63 = ~ T64;
  assign T64 = 4'h0 - T155;
  assign T155 = {3'h0, T65};
  assign T65 = T71 & T66;
  assign T66 = T68 | T67;
  assign T67 = 3'h2 == io_inner_release_bits_r_type;
  assign T68 = T70 | T69;
  assign T69 = 3'h1 == io_inner_release_bits_r_type;
  assign T70 = 3'h0 == io_inner_release_bits_r_type;
  assign T71 = io_inner_release_ready & io_inner_release_valid;
  assign T72 = T75 | T73;
  assign T73 = ~ T74;
  assign T74 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T75 = ~ T76;
  assign T76 = 4'h0 - T156;
  assign T156 = {3'h0, T77};
  assign T77 = T83 & T78;
  assign T78 = T80 | T79;
  assign T79 = 3'h2 == io_inner_release_bits_r_type;
  assign T80 = T82 | T81;
  assign T81 = 3'h1 == io_inner_release_bits_r_type;
  assign T82 = 3'h0 == io_inner_release_bits_r_type;
  assign T83 = io_inner_release_ready & io_inner_release_valid;
  assign T84 = T10 & T85;
  assign T85 = T87 | T86;
  assign T86 = 3'h2 == io_inner_release_bits_r_type;
  assign T87 = T89 | T88;
  assign T88 = 3'h1 == io_inner_release_bits_r_type;
  assign T89 = 3'h0 == io_inner_release_bits_r_type;
  assign T90 = T10 & T91;
  assign T91 = T85 ^ 1'h1;
  assign T92 = state == 1'h1;
  assign io_has_acquire_match = 1'h0;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = T93;
  assign T93 = T94 & io_inner_grant_ready;
  assign T94 = state == 1'h1;
  assign io_outer_acquire_bits_data = T95;
  assign T95 = T96;
  assign T96 = T117 ? T109 : T97;
  assign T97 = T107 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T98 = T99 ? io_inner_release_bits_data : xact_data_buffer_0;
  assign T99 = T103 & T100;
  assign T100 = T101[1'h0];
  assign T101 = 1'h1 << T102;
  assign T102 = io_inner_release_bits_addr_beat;
  assign T103 = io_inner_release_ready & io_inner_release_valid;
  assign T104 = T105 ? io_inner_release_bits_data : xact_data_buffer_1;
  assign T105 = T103 & T106;
  assign T106 = T101[1'h1];
  assign T107 = T108[1'h0];
  assign T108 = T157;
  assign T157 = T162 ? 1'h0 : T158;
  assign T158 = T161 ? 1'h1 : T159;
  assign T159 = T160 ? 2'h2 : 2'h3;
  assign T160 = pending_writes[2'h2];
  assign T161 = pending_writes[1'h1];
  assign T162 = pending_writes[1'h0];
  assign T109 = T116 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T110 = T111 ? io_inner_release_bits_data : xact_data_buffer_2;
  assign T111 = T103 & T112;
  assign T112 = T101[2'h2];
  assign T113 = T114 ? io_inner_release_bits_data : xact_data_buffer_3;
  assign T114 = T103 & T115;
  assign T115 = T101[2'h3];
  assign T116 = T108[1'h0];
  assign T117 = T108[1'h1];
  assign io_outer_acquire_bits_union = T118;
  assign T118 = T119;
  assign T119 = {T120, 1'h1};
  assign T120 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T121;
  assign T121 = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T122;
  assign T122 = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T123;
  assign T123 = T157;
  assign io_outer_acquire_bits_client_xact_id = T163;
  assign T163 = T124[2'h3:1'h0];
  assign T124 = 6'h0;
  assign io_outer_acquire_bits_addr_block = T125;
  assign T125 = xact_addr_block;
  assign T126 = T10 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign io_outer_acquire_valid = T127;
  assign T127 = T129 & T128;
  assign T128 = pending_writes != 4'h0;
  assign T129 = state == 1'h1;
  assign io_inner_release_ready = T130;
  assign T130 = T132 | T131;
  assign T131 = pending_irels != 4'h0;
  assign T132 = T133 & io_inner_release_bits_voluntary;
  assign T133 = state == 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_grant_bits_client_id = T134;
  assign T134 = xact_client_id;
  assign T135 = T10 ? io_inner_release_bits_client_id : xact_client_id;
  assign io_inner_grant_bits_data = T136;
  assign T136 = 4'h0;
  assign io_inner_grant_bits_g_type = T137;
  assign T137 = 4'h0;
  assign io_inner_grant_bits_is_builtin_type = T138;
  assign T138 = 1'h1;
  assign io_inner_grant_bits_manager_xact_id = T139;
  assign T139 = 4'h0;
  assign io_inner_grant_bits_client_xact_id = T140;
  assign T140 = xact_client_xact_id;
  assign T141 = T10 ? io_inner_release_bits_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T142;
  assign T142 = 2'h0;
  assign io_inner_grant_valid = T143;
  assign T143 = T144 & io_outer_grant_valid;
  assign T144 = T146 & T145;
  assign T145 = pending_irels == 4'h0;
  assign T146 = T147 & pending_ignt;
  assign T147 = state == 1'h1;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "VoluntaryReleaseTracker accepted Release that wasn't voluntary!");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 1'h0;
    end else if(T13) begin
      state <= 1'h0;
    end else if(T10) begin
      state <= 1'h1;
    end
    if(reset) begin
      pending_ignt <= 1'h0;
    end else if(T10) begin
      pending_ignt <= 1'h1;
    end else if(T17) begin
      pending_ignt <= 1'h0;
    end
    if(reset) begin
      pending_writes <= 4'h0;
    end else if(T10) begin
      pending_writes <= T46;
    end else begin
      pending_writes <= T21;
    end
    if(reset) begin
      pending_irels <= 4'h0;
    end else if(T90) begin
      pending_irels <= 4'h0;
    end else if(T84) begin
      pending_irels <= T72;
    end else begin
      pending_irels <= T59;
    end
    if(T99) begin
      xact_data_buffer_0 <= io_inner_release_bits_data;
    end
    if(T105) begin
      xact_data_buffer_1 <= io_inner_release_bits_data;
    end
    if(T111) begin
      xact_data_buffer_2 <= io_inner_release_bits_data;
    end
    if(T114) begin
      xact_data_buffer_3 <= io_inner_release_bits_data;
    end
    if(T10) begin
      xact_addr_block <= io_inner_release_bits_addr_block;
    end
    if(T10) begin
      xact_client_id <= io_inner_release_bits_client_id;
    end
    if(T10) begin
      xact_client_xact_id <= io_inner_release_bits_client_xact_id;
    end
  end
endmodule

module BroadcastAcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h1;
  assign oacq_read_beat_client_xact_id = 4'h1;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h1;
  assign oacq_write_beat_client_xact_id = 4'h1;
  assign oacq_probe_client_xact_id = 4'h1;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h1;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h2;
  assign oacq_read_beat_client_xact_id = 4'h2;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h2;
  assign oacq_write_beat_client_xact_id = 4'h2;
  assign oacq_probe_client_xact_id = 4'h2;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h2;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h3;
  assign oacq_read_beat_client_xact_id = 4'h3;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h3;
  assign oacq_write_beat_client_xact_id = 4'h3;
  assign oacq_probe_client_xact_id = 4'h3;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h3;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h4;
  assign oacq_read_beat_client_xact_id = 4'h4;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h4;
  assign oacq_write_beat_client_xact_id = 4'h4;
  assign oacq_probe_client_xact_id = 4'h4;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h4;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h5;
  assign oacq_read_beat_client_xact_id = 4'h5;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h5;
  assign oacq_write_beat_client_xact_id = 4'h5;
  assign oacq_probe_client_xact_id = 4'h5;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h5;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h6;
  assign oacq_read_beat_client_xact_id = 4'h6;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h6;
  assign oacq_write_beat_client_xact_id = 4'h6;
  assign oacq_probe_client_xact_id = 4'h6;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h6;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module BroadcastAcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T477;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T478;
  wire[2:0] T25;
  wire[2:0] T479;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T480;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T481;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T482;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T483;
  wire[2:0] T484;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T485;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T486;
  wire T88;
  wire[2:0] T487;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T488;
  wire T92;
  wire T93;
  wire[2:0] T489;
  wire T94;
  wire[2:0] T490;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [25:0] xact_addr_block;
  wire[25:0] T108;
  wire T109;
  wire T110;
  wire oacq_data_done;
  wire T111;
  wire T112;
  wire T113;
  reg [1:0] R114;
  wire[1:0] T491;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire[2:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire ignt_data_done;
  wire T137;
  wire T138;
  wire T139;
  reg [1:0] R140;
  wire[1:0] T492;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  reg [5:0] xact_client_xact_id;
  wire[5:0] T163;
  wire T164;
  wire T165;
  wire T166;
  reg  collect_iacq_data;
  wire T493;
  wire T167;
  wire T168;
  wire T169;
  wire iacq_data_done;
  wire T170;
  wire T171;
  wire T172;
  reg [1:0] R173;
  wire[1:0] T494;
  wire[1:0] T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg  T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg [1:0] xact_client_id;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg  pending_ognt_ack;
  wire T495;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T224;
  wire[3:0] T225;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T226;
  wire[3:0] T227;
  wire T228;
  wire T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T237;
  wire[3:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T245;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T246;
  wire[3:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T252;
  wire[3:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[3:0] oacq_write_beat_data;
  wire T260;
  wire[3:0] oacq_probe_data;
  wire T261;
  wire[16:0] T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T496;
  wire[12:0] T265;
  wire[6:0] T266;
  wire[2:0] T267;
  reg [16:0] xact_union;
  wire[16:0] T268;
  wire[3:0] T269;
  wire[16:0] T270;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T271;
  wire[15:0] T272;
  wire[15:0] T273;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[15:0] T284;
  wire[15:0] T285;
  wire[7:0] T286;
  wire[7:0] T497;
  wire T287;
  wire[1:0] T288;
  wire T289;
  wire[3:0] T290;
  wire[7:0] T291;
  wire[7:0] T498;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[15:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire[15:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[7:0] T499;
  wire T310;
  wire[1:0] T311;
  wire T312;
  wire[3:0] T313;
  wire[7:0] T314;
  wire[7:0] T500;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[3:0] T320;
  wire[1:0] T321;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T322;
  wire[15:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[15:0] T330;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T331;
  wire[15:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T337;
  wire[15:0] T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T345;
  wire[15:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[15:0] T354;
  wire[15:0] T355;
  wire[7:0] T356;
  wire[7:0] T501;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[7:0] T361;
  wire[7:0] T502;
  wire T362;
  wire T363;
  wire T364;
  wire[16:0] oacq_probe_union;
  wire[16:0] T365;
  wire[15:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T370;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T371;
  wire T372;
  wire T373;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T374;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] oacq_read_block_client_xact_id;
  wire[3:0] oacq_read_beat_client_xact_id;
  wire[3:0] T383;
  wire[3:0] oacq_write_block_client_xact_id;
  wire[3:0] oacq_write_beat_client_xact_id;
  wire[3:0] oacq_probe_client_xact_id;
  wire[25:0] T384;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T387;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg [3:0] iacq_data_valid;
  wire[3:0] T503;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[3:0] T504;
  wire T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T505;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[25:0] T447;
  wire T448;
  wire T449;
  reg  pending_probes;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T421;
  wire[3:0] T422;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[1:0] T510;
  wire T426;
  wire[1:0] T450;
  wire[3:0] T451;
  wire[3:0] T452;
  wire[3:0] T511;
  wire[2:0] T453;
  wire[2:0] T512;
  wire[1:0] T454;
  wire T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire[2:0] T458;
  wire[2:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[5:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    xact_addr_block = {1{$random}};
    R114 = {1{$random}};
    R140 = {1{$random}};
    T158 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R173 = {1{$random}};
    T182 = 1'b0;
    xact_client_id = {1{$random}};
    T192 = 1'b0;
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T477 = reset ? 3'h0 : T11;
  assign T11 = T156 ? 3'h0 : T12;
  assign T12 = T154 ? T150 : T13;
  assign T13 = T136 ? T132 : T14;
  assign T14 = T129 ? 3'h5 : T15;
  assign T15 = T127 ? T126 : T16;
  assign T16 = T124 ? T122 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T478;
  assign T478 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T479;
  assign T479 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T480;
  assign T480 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T481 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T481 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T482 & T59;
  assign T59 = ~ T56;
  assign T482 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T110 & T79;
  assign T79 = release_count == 1'h1;
  assign T483 = T484[1'h0];
  assign T484 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T490 : T81;
  assign T81 = T110 ? T489 : T82;
  assign T82 = T93 ? T83 : T485;
  assign T485 = {2'h0, release_count};
  assign T83 = T487 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T486 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3];
  assign T486 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2];
  assign T487 = {1'h0, T89};
  assign T89 = T488 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1];
  assign T488 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0];
  assign T93 = T61 & T52;
  assign T489 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T490 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T109 & T104;
  assign T104 = io_inner_release_valid & T105;
  assign T105 = T107 & T106;
  assign T106 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T107 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T108 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign T109 = 3'h1 == state;
  assign T110 = T120 & oacq_data_done;
  assign oacq_data_done = T118 ? T112 : T111;
  assign T111 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T112 = T117 & T113;
  assign T113 = R114 == 2'h3;
  assign T491 = reset ? 2'h0 : T115;
  assign T115 = T117 ? T116 : R114;
  assign T116 = R114 + 2'h1;
  assign T117 = T111 & T118;
  assign T118 = io_outer_acquire_bits_is_builtin_type & T119;
  assign T119 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T120 = T121 & io_outer_acquire_ready;
  assign T121 = T103 & T98;
  assign T122 = pending_outer_write ? 3'h3 : T123;
  assign T123 = pending_outer_read ? 3'h2 : 3'h4;
  assign T124 = T96 & T125;
  assign T125 = release_count == 1'h1;
  assign T126 = pending_outer_read ? 3'h2 : 3'h5;
  assign T127 = T128 & oacq_data_done;
  assign T128 = 3'h3 == state;
  assign T129 = T131 & T130;
  assign T130 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T131 = 3'h2 == state;
  assign T132 = T133 ? 3'h6 : 3'h0;
  assign T133 = T134 ^ 1'h1;
  assign T134 = io_inner_grant_bits_is_builtin_type & T135;
  assign T135 = io_inner_grant_bits_g_type == 4'h0;
  assign T136 = T149 & ignt_data_done;
  assign ignt_data_done = T144 ? T138 : T137;
  assign T137 = io_inner_grant_ready & io_inner_grant_valid;
  assign T138 = T143 & T139;
  assign T139 = R140 == 2'h3;
  assign T492 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : R140;
  assign T142 = R140 + 2'h1;
  assign T143 = T137 & T144;
  assign T144 = io_inner_grant_bits_is_builtin_type ? T148 : T145;
  assign T145 = T147 | T146;
  assign T146 = 4'h1 == io_inner_grant_bits_g_type;
  assign T147 = 4'h0 == io_inner_grant_bits_g_type;
  assign T148 = 4'h5 == io_inner_grant_bits_g_type;
  assign T149 = 3'h5 == state;
  assign T150 = T151 ? 3'h6 : 3'h0;
  assign T151 = T152 ^ 1'h1;
  assign T152 = io_inner_grant_bits_is_builtin_type & T153;
  assign T153 = io_inner_grant_bits_g_type == 4'h0;
  assign T154 = T155 & io_inner_grant_ready;
  assign T155 = 3'h4 == state;
  assign T156 = T157 & io_inner_finish_valid;
  assign T157 = 3'h6 == state;
  assign T159 = T160 | reset;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T164 & T162;
  assign T162 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T163 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T164 = T166 & T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T181 & collect_iacq_data;
  assign T493 = reset ? 1'h0 : T167;
  assign T167 = T61 ? T179 : T168;
  assign T168 = T169 ? 1'h0 : collect_iacq_data;
  assign T169 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T177 ? T171 : T170;
  assign T170 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T171 = T176 & T172;
  assign T172 = R173 == 2'h3;
  assign T494 = reset ? 2'h0 : T174;
  assign T174 = T176 ? T175 : R173;
  assign T175 = R173 + 2'h1;
  assign T176 = T170 & T177;
  assign T177 = io_inner_acquire_bits_is_builtin_type & T178;
  assign T178 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T179 = io_inner_acquire_bits_is_builtin_type & T180;
  assign T180 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T188 & T186;
  assign T186 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T187 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T188 = T190 & T189;
  assign T189 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T190 = T191 & collect_iacq_data;
  assign T191 = state != 3'h0;
  assign T193 = T194 | reset;
  assign T194 = T195 ^ 1'h1;
  assign T195 = T201 & T196;
  assign T196 = T198 | T197;
  assign T197 = 3'h6 == xact_a_type;
  assign T198 = T200 | T199;
  assign T199 = 3'h5 == xact_a_type;
  assign T200 = 3'h4 == xact_a_type;
  assign T201 = T202 & xact_is_builtin_type;
  assign T202 = state != 3'h0;
  assign io_has_acquire_match = T203;
  assign T203 = T204 & collect_iacq_data;
  assign T204 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T205;
  assign T205 = T207 & T206;
  assign T206 = collect_iacq_data ^ 1'h1;
  assign T207 = T209 & T208;
  assign T208 = state != 3'h0;
  assign T209 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T210;
  assign T210 = T149 ? io_inner_grant_ready : pending_ognt_ack;
  assign T495 = reset ? 1'h0 : T211;
  assign T211 = T127 ? 1'h1 : T212;
  assign T212 = T110 ? 1'h1 : T213;
  assign T213 = T214 ? 1'h0 : pending_ognt_ack;
  assign T214 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T215;
  assign T215 = T261 ? oacq_probe_data : T216;
  assign T216 = T260 ? T223 : T217;
  assign T217 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T218;
  assign T218 = T220 | T219;
  assign T219 = 3'h4 == xact_a_type;
  assign T220 = T222 | T221;
  assign T221 = 3'h0 == xact_a_type;
  assign T222 = 3'h2 == xact_a_type;
  assign T223 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T224;
  assign T224 = T259 ? T245 : T225;
  assign T225 = T243 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T226 = T233 ? io_inner_acquire_bits_data : T227;
  assign T227 = T228 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T228 = T232 & T229;
  assign T229 = T230[1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = io_inner_acquire_bits_addr_beat;
  assign T232 = collect_iacq_data & io_inner_acquire_valid;
  assign T233 = T61 & T234;
  assign T234 = T235[1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = 2'h0;
  assign T237 = T241 ? io_inner_acquire_bits_data : T238;
  assign T238 = T239 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T239 = T232 & T240;
  assign T240 = T230[1'h1];
  assign T241 = T61 & T242;
  assign T242 = T235[1'h1];
  assign T243 = T244[1'h0];
  assign T244 = oacq_data_cnt;
  assign oacq_data_cnt = T118 ? R114 : 2'h0;
  assign T245 = T258 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T246 = T250 ? io_inner_acquire_bits_data : T247;
  assign T247 = T248 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T248 = T232 & T249;
  assign T249 = T230[2'h2];
  assign T250 = T61 & T251;
  assign T251 = T235[2'h2];
  assign T252 = T256 ? io_inner_acquire_bits_data : T253;
  assign T253 = T254 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T254 = T232 & T255;
  assign T255 = T230[2'h3];
  assign T256 = T61 & T257;
  assign T257 = T235[2'h3];
  assign T258 = T244[1'h0];
  assign T259 = T244[1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T260 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T261 = state == 3'h1;
  assign io_outer_acquire_bits_union = T262;
  assign T262 = T261 ? oacq_probe_union : T263;
  assign T263 = T260 ? T270 : T264;
  assign T264 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T496;
  assign T496 = {4'h0, T265};
  assign T265 = {T266, 6'h0};
  assign T266 = {T269, T267};
  assign T267 = xact_union[4'h8:3'h6];
  assign T268 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T269 = xact_union[4'hc:4'h9];
  assign T270 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T271;
  assign T271 = {T272, 1'h1};
  assign T272 = T344 ? T330 : T273;
  assign T273 = T328 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T274 = T318 ? T299 : T275;
  assign T275 = T295 ? T276 : xact_wmask_buffer_0;
  assign T276 = T293 ? T284 : T277;
  assign T277 = T279 ? T278 : 16'h0;
  assign T278 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T279 = T282 | T280;
  assign T280 = io_inner_acquire_bits_is_builtin_type & T281;
  assign T281 = io_inner_acquire_bits_a_type == 3'h2;
  assign T282 = io_inner_acquire_bits_is_builtin_type & T283;
  assign T283 = io_inner_acquire_bits_a_type == 3'h3;
  assign T284 = T285;
  assign T285 = {T291, T286};
  assign T286 = 8'h0 - T497;
  assign T497 = {7'h0, T287};
  assign T287 = T288[1'h0];
  assign T288 = 1'h1 << T289;
  assign T289 = T290[2'h3];
  assign T290 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T291 = 8'h0 - T498;
  assign T498 = {7'h0, T292};
  assign T292 = T288[1'h1];
  assign T293 = io_inner_acquire_bits_is_builtin_type & T294;
  assign T294 = io_inner_acquire_bits_a_type == 3'h4;
  assign T295 = T232 & T296;
  assign T296 = T297[1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = io_inner_acquire_bits_addr_beat;
  assign T299 = T316 ? T307 : T300;
  assign T300 = T302 ? T301 : 16'h0;
  assign T301 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T302 = T305 | T303;
  assign T303 = io_inner_acquire_bits_is_builtin_type & T304;
  assign T304 = io_inner_acquire_bits_a_type == 3'h2;
  assign T305 = io_inner_acquire_bits_is_builtin_type & T306;
  assign T306 = io_inner_acquire_bits_a_type == 3'h3;
  assign T307 = T308;
  assign T308 = {T314, T309};
  assign T309 = 8'h0 - T499;
  assign T499 = {7'h0, T310};
  assign T310 = T311[1'h0];
  assign T311 = 1'h1 << T312;
  assign T312 = T313[2'h3];
  assign T313 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T314 = 8'h0 - T500;
  assign T500 = {7'h0, T315};
  assign T315 = T311[1'h1];
  assign T316 = io_inner_acquire_bits_is_builtin_type & T317;
  assign T317 = io_inner_acquire_bits_a_type == 3'h4;
  assign T318 = T61 & T319;
  assign T319 = T320[1'h0];
  assign T320 = 1'h1 << T321;
  assign T321 = 2'h0;
  assign T322 = T326 ? T299 : T323;
  assign T323 = T324 ? T276 : xact_wmask_buffer_1;
  assign T324 = T232 & T325;
  assign T325 = T297[1'h1];
  assign T326 = T61 & T327;
  assign T327 = T320[1'h1];
  assign T328 = T329[1'h0];
  assign T329 = oacq_data_cnt;
  assign T330 = T343 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T331 = T335 ? T299 : T332;
  assign T332 = T333 ? T276 : xact_wmask_buffer_2;
  assign T333 = T232 & T334;
  assign T334 = T297[2'h2];
  assign T335 = T61 & T336;
  assign T336 = T320[2'h2];
  assign T337 = T341 ? T299 : T338;
  assign T338 = T339 ? T276 : xact_wmask_buffer_3;
  assign T339 = T232 & T340;
  assign T340 = T297[2'h3];
  assign T341 = T61 & T342;
  assign T342 = T320[2'h3];
  assign T343 = T329[1'h0];
  assign T344 = T329[1'h1];
  assign oacq_write_beat_union = T345;
  assign T345 = {T346, 1'h1};
  assign T346 = T363 ? T354 : T347;
  assign T347 = T349 ? T348 : 16'h0;
  assign T348 = xact_union[5'h10:1'h1];
  assign T349 = T352 | T350;
  assign T350 = xact_is_builtin_type & T351;
  assign T351 = xact_a_type == 3'h2;
  assign T352 = xact_is_builtin_type & T353;
  assign T353 = xact_a_type == 3'h3;
  assign T354 = T355;
  assign T355 = {T361, T356};
  assign T356 = 8'h0 - T501;
  assign T501 = {7'h0, T357};
  assign T357 = T358[1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = T360[2'h3];
  assign T360 = xact_union[4'hc:4'h9];
  assign T361 = 8'h0 - T502;
  assign T502 = {7'h0, T362};
  assign T362 = T358[1'h1];
  assign T363 = xact_is_builtin_type & T364;
  assign T364 = xact_a_type == 3'h4;
  assign oacq_probe_union = T365;
  assign T365 = {T366, 1'h1};
  assign T366 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T367;
  assign T367 = T261 ? oacq_probe_a_type : T368;
  assign T368 = T260 ? T370 : T369;
  assign T369 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T370 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T371;
  assign T371 = T261 ? oacq_probe_is_builtin_type : T372;
  assign T372 = T260 ? T374 : T373;
  assign T373 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T374 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T375;
  assign T375 = T261 ? oacq_probe_addr_beat : T376;
  assign T376 = T260 ? T379 : T377;
  assign T377 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T378 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T379 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T380;
  assign T380 = T261 ? oacq_probe_client_xact_id : T381;
  assign T381 = T260 ? T383 : T382;
  assign T382 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 4'h7;
  assign oacq_read_beat_client_xact_id = 4'h7;
  assign T383 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 4'h7;
  assign oacq_write_beat_client_xact_id = 4'h7;
  assign oacq_probe_client_xact_id = 4'h7;
  assign io_outer_acquire_bits_addr_block = T384;
  assign T384 = T261 ? oacq_probe_addr_block : T385;
  assign T385 = T260 ? T387 : T386;
  assign T386 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T387 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T388;
  assign T388 = T131 ? T410 : T389;
  assign T389 = T128 ? T390 : T121;
  assign T390 = T409 & T391;
  assign T391 = T408 | T392;
  assign T392 = iacq_data_valid[oacq_data_cnt];
  assign T503 = reset ? 4'h0 : T393;
  assign T393 = T61 ? T401 : T394;
  assign T394 = T232 ? T395 : iacq_data_valid;
  assign T395 = T399 | T396;
  assign T396 = T504 & T397;
  assign T397 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T504 = T398 ? 4'hf : 4'h0;
  assign T398 = 1'h1;
  assign T399 = iacq_data_valid & T400;
  assign T400 = ~ T397;
  assign T401 = T402 << io_inner_acquire_bits_addr_beat;
  assign T402 = io_inner_acquire_bits_is_builtin_type & T403;
  assign T403 = T405 | T404;
  assign T404 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T405 = T407 | T406;
  assign T406 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T407 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T408 = collect_iacq_data ^ 1'h1;
  assign T409 = pending_ognt_ack ^ 1'h1;
  assign T410 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T411;
  assign T411 = T109 ? T412 : 1'h0;
  assign T412 = T413 & T105;
  assign T413 = T414 | io_outer_acquire_ready;
  assign T414 = T415 ^ 1'h1;
  assign T415 = T417 | T416;
  assign T416 = 3'h2 == io_inner_release_bits_r_type;
  assign T417 = T419 | T418;
  assign T418 = 3'h1 == io_inner_release_bits_r_type;
  assign T419 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T420;
  assign T420 = T505;
  assign T505 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T427;
  assign T427 = T428;
  assign T428 = xact_is_builtin_type ? T433 : T429;
  assign T429 = T432 ? 2'h1 : T430;
  assign T430 = T431 ? 2'h0 : 2'h2;
  assign T431 = xact_a_type == 3'h1;
  assign T432 = xact_a_type == 3'h0;
  assign T433 = T446 ? 2'h2 : T434;
  assign T434 = T445 ? 2'h0 : T435;
  assign T435 = T444 ? 2'h2 : T436;
  assign T436 = T443 ? 2'h0 : T437;
  assign T437 = T442 ? 2'h2 : T438;
  assign T438 = T441 ? 2'h0 : T439;
  assign T439 = T440 ? 2'h0 : 2'h2;
  assign T440 = xact_a_type == 3'h4;
  assign T441 = xact_a_type == 3'h6;
  assign T442 = xact_a_type == 3'h5;
  assign T443 = xact_a_type == 3'h2;
  assign T444 = xact_a_type == 3'h0;
  assign T445 = xact_a_type == 3'h3;
  assign T446 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T447;
  assign T447 = xact_addr_block;
  assign io_inner_probe_valid = T448;
  assign T448 = T109 ? T449 : 1'h0;
  assign T449 = pending_probes != 1'h0;
  assign T506 = T507[1'h0];
  assign T507 = reset ? 4'h0 : T421;
  assign T421 = T426 ? T509 : T422;
  assign T422 = T93 ? mask_incoherent : T508;
  assign T508 = {3'h0, pending_probes};
  assign T509 = {2'h0, T423};
  assign T423 = T510 & T424;
  assign T424 = ~ T425;
  assign T425 = 1'h1 << 1'h0;
  assign T510 = {1'h0, pending_probes};
  assign T426 = T109 & io_inner_probe_ready;
  assign io_inner_finish_ready = T157;
  assign io_inner_grant_bits_client_id = T450;
  assign T450 = xact_client_id;
  assign io_inner_grant_bits_data = T451;
  assign T451 = 4'h0;
  assign io_inner_grant_bits_g_type = T452;
  assign T452 = T511;
  assign T511 = {1'h0, T453};
  assign T453 = xact_is_builtin_type ? T456 : T512;
  assign T512 = {1'h0, T454};
  assign T454 = T455 ? 2'h0 : 2'h1;
  assign T455 = xact_a_type == 3'h0;
  assign T456 = T469 ? 3'h4 : T457;
  assign T457 = T468 ? 3'h5 : T458;
  assign T458 = T467 ? 3'h3 : T459;
  assign T459 = T466 ? 3'h3 : T460;
  assign T460 = T465 ? 3'h4 : T461;
  assign T461 = T464 ? 3'h1 : T462;
  assign T462 = T463 ? 3'h1 : 3'h3;
  assign T463 = xact_a_type == 3'h6;
  assign T464 = xact_a_type == 3'h5;
  assign T465 = xact_a_type == 3'h4;
  assign T466 = xact_a_type == 3'h3;
  assign T467 = xact_a_type == 3'h2;
  assign T468 = xact_a_type == 3'h1;
  assign T469 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T470;
  assign T470 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T471;
  assign T471 = 4'h7;
  assign io_inner_grant_bits_client_xact_id = T472;
  assign T472 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T473;
  assign T473 = 2'h0;
  assign io_inner_grant_valid = T474;
  assign T474 = T155 ? 1'h1 : T475;
  assign T475 = T149 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T476;
  assign T476 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T192 <= 1'b1;
  if(!T193 && T192 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T158 <= 1'b1;
  if(!T159 && T158 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T156) begin
      state <= 3'h0;
    end else if(T154) begin
      state <= T150;
    end else if(T136) begin
      state <= T132;
    end else if(T129) begin
      state <= 3'h5;
    end else if(T127) begin
      state <= T126;
    end else if(T124) begin
      state <= T122;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T483;
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      R114 <= 2'h0;
    end else if(T117) begin
      R114 <= T116;
    end
    if(reset) begin
      R140 <= 2'h0;
    end else if(T143) begin
      R140 <= T142;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T179;
    end else if(T169) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R173 <= 2'h0;
    end else if(T176) begin
      R173 <= T175;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T127) begin
      pending_ognt_ack <= 1'h1;
    end else if(T110) begin
      pending_ognt_ack <= 1'h1;
    end else if(T214) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T233) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T228) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T241) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T239) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T250) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T248) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T256) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T254) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T318) begin
      xact_wmask_buffer_0 <= T299;
    end else if(T295) begin
      xact_wmask_buffer_0 <= T276;
    end
    if(T326) begin
      xact_wmask_buffer_1 <= T299;
    end else if(T324) begin
      xact_wmask_buffer_1 <= T276;
    end
    if(T335) begin
      xact_wmask_buffer_2 <= T299;
    end else if(T333) begin
      xact_wmask_buffer_2 <= T276;
    end
    if(T341) begin
      xact_wmask_buffer_3 <= T299;
    end else if(T339) begin
      xact_wmask_buffer_3 <= T276;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T401;
    end else if(T232) begin
      iacq_data_valid <= T395;
    end
    pending_probes <= T506;
  end
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_addr_beat,
    input [5:0] io_in_7_bits_client_xact_id,
    input [3:0] io_in_7_bits_manager_xact_id,
    input  io_in_7_bits_is_builtin_type,
    input [3:0] io_in_7_bits_g_type,
    input [127:0] io_in_7_bits_data,
    input [1:0] io_in_7_bits_client_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_addr_beat,
    input [5:0] io_in_6_bits_client_xact_id,
    input [3:0] io_in_6_bits_manager_xact_id,
    input  io_in_6_bits_is_builtin_type,
    input [3:0] io_in_6_bits_g_type,
    input [127:0] io_in_6_bits_data,
    input [1:0] io_in_6_bits_client_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_addr_beat,
    input [5:0] io_in_5_bits_client_xact_id,
    input [3:0] io_in_5_bits_manager_xact_id,
    input  io_in_5_bits_is_builtin_type,
    input [3:0] io_in_5_bits_g_type,
    input [127:0] io_in_5_bits_data,
    input [1:0] io_in_5_bits_client_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_addr_beat,
    input [5:0] io_in_4_bits_client_xact_id,
    input [3:0] io_in_4_bits_manager_xact_id,
    input  io_in_4_bits_is_builtin_type,
    input [3:0] io_in_4_bits_g_type,
    input [127:0] io_in_4_bits_data,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_addr_beat,
    input [5:0] io_in_3_bits_client_xact_id,
    input [3:0] io_in_3_bits_manager_xact_id,
    input  io_in_3_bits_is_builtin_type,
    input [3:0] io_in_3_bits_g_type,
    input [127:0] io_in_3_bits_data,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_addr_beat,
    input [5:0] io_in_2_bits_client_xact_id,
    input [3:0] io_in_2_bits_manager_xact_id,
    input  io_in_2_bits_is_builtin_type,
    input [3:0] io_in_2_bits_g_type,
    input [127:0] io_in_2_bits_data,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [5:0] io_in_1_bits_client_xact_id,
    input [3:0] io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [127:0] io_in_1_bits_data,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [5:0] io_in_0_bits_client_xact_id,
    input [3:0] io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [127:0] io_in_0_bits_data,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[5:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T359;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T360;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  reg  locked;
  wire T361;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  reg [1:0] R59;
  wire[1:0] T362;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire T66;
  wire[2:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire T73;
  wire[1:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire[127:0] T78;
  wire[127:0] T79;
  wire[127:0] T80;
  wire T81;
  wire[127:0] T82;
  wire T83;
  wire T84;
  wire[127:0] T85;
  wire[127:0] T86;
  wire T87;
  wire[127:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[3:0] T94;
  wire T95;
  wire[3:0] T96;
  wire T97;
  wire T98;
  wire[3:0] T99;
  wire[3:0] T100;
  wire T101;
  wire[3:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire T123;
  wire[3:0] T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[5:0] T134;
  wire[5:0] T135;
  wire[5:0] T136;
  wire T137;
  wire[5:0] T138;
  wire T139;
  wire T140;
  wire[5:0] T141;
  wire[5:0] T142;
  wire T143;
  wire[5:0] T144;
  wire T145;
  wire T146;
  wire T147;
  wire[1:0] T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire T151;
  wire[1:0] T152;
  wire T153;
  wire T154;
  wire[1:0] T155;
  wire[1:0] T156;
  wire T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R59 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T359 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T360 = reset ? 3'h7 : T30;
  assign T30 = T45 ? T31 : lockIdx;
  assign T31 = T44 ? 3'h0 : T32;
  assign T32 = T43 ? 3'h1 : T33;
  assign T33 = T42 ? 3'h2 : T34;
  assign T34 = T41 ? 3'h3 : T35;
  assign T35 = T40 ? 3'h4 : T36;
  assign T36 = T39 ? 3'h5 : T37;
  assign T37 = T38 ? 3'h6 : 3'h7;
  assign T38 = io_in_6_ready & io_in_6_valid;
  assign T39 = io_in_5_ready & io_in_5_valid;
  assign T40 = io_in_4_ready & io_in_4_valid;
  assign T41 = io_in_3_ready & io_in_3_valid;
  assign T42 = io_in_2_ready & io_in_2_valid;
  assign T43 = io_in_1_ready & io_in_1_valid;
  assign T44 = io_in_0_ready & io_in_0_valid;
  assign T45 = T47 & T46;
  assign T46 = locked ^ 1'h1;
  assign T47 = T53 & T48;
  assign T48 = io_out_bits_is_builtin_type ? T52 : T49;
  assign T49 = T51 | T50;
  assign T50 = 4'h1 == io_out_bits_g_type;
  assign T51 = 4'h0 == io_out_bits_g_type;
  assign T52 = 4'h5 == io_out_bits_g_type;
  assign T53 = io_out_valid & io_out_ready;
  assign T361 = reset ? 1'h0 : T54;
  assign T54 = T61 ? 1'h0 : T55;
  assign T55 = T47 ? T56 : locked;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T58 == 2'h0;
  assign T58 = R59 + 2'h1;
  assign T362 = reset ? 2'h0 : T60;
  assign T60 = T47 ? T58 : R59;
  assign T61 = T53 & T62;
  assign T62 = T48 ^ 1'h1;
  assign io_out_bits_client_id = T63;
  assign T63 = T77 ? T71 : T64;
  assign T64 = T70 ? T68 : T65;
  assign T65 = T66 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T66 = T67[1'h0];
  assign T67 = chosen;
  assign T68 = T69 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T69 = T67[1'h0];
  assign T70 = T67[1'h1];
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? io_in_5_bits_client_id : io_in_4_bits_client_id;
  assign T73 = T67[1'h0];
  assign T74 = T75 ? io_in_7_bits_client_id : io_in_6_bits_client_id;
  assign T75 = T67[1'h0];
  assign T76 = T67[1'h1];
  assign T77 = T67[2'h2];
  assign io_out_bits_data = T78;
  assign T78 = T91 ? T85 : T79;
  assign T79 = T84 ? T82 : T80;
  assign T80 = T81 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T81 = T67[1'h0];
  assign T82 = T83 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T83 = T67[1'h0];
  assign T84 = T67[1'h1];
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? io_in_5_bits_data : io_in_4_bits_data;
  assign T87 = T67[1'h0];
  assign T88 = T89 ? io_in_7_bits_data : io_in_6_bits_data;
  assign T89 = T67[1'h0];
  assign T90 = T67[1'h1];
  assign T91 = T67[2'h2];
  assign io_out_bits_g_type = T92;
  assign T92 = T105 ? T99 : T93;
  assign T93 = T98 ? T96 : T94;
  assign T94 = T95 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign T95 = T67[1'h0];
  assign T96 = T97 ? io_in_3_bits_g_type : io_in_2_bits_g_type;
  assign T97 = T67[1'h0];
  assign T98 = T67[1'h1];
  assign T99 = T104 ? T102 : T100;
  assign T100 = T101 ? io_in_5_bits_g_type : io_in_4_bits_g_type;
  assign T101 = T67[1'h0];
  assign T102 = T103 ? io_in_7_bits_g_type : io_in_6_bits_g_type;
  assign T103 = T67[1'h0];
  assign T104 = T67[1'h1];
  assign T105 = T67[2'h2];
  assign io_out_bits_is_builtin_type = T106;
  assign T106 = T119 ? T113 : T107;
  assign T107 = T112 ? T110 : T108;
  assign T108 = T109 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T109 = T67[1'h0];
  assign T110 = T111 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T111 = T67[1'h0];
  assign T112 = T67[1'h1];
  assign T113 = T118 ? T116 : T114;
  assign T114 = T115 ? io_in_5_bits_is_builtin_type : io_in_4_bits_is_builtin_type;
  assign T115 = T67[1'h0];
  assign T116 = T117 ? io_in_7_bits_is_builtin_type : io_in_6_bits_is_builtin_type;
  assign T117 = T67[1'h0];
  assign T118 = T67[1'h1];
  assign T119 = T67[2'h2];
  assign io_out_bits_manager_xact_id = T120;
  assign T120 = T133 ? T127 : T121;
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign T123 = T67[1'h0];
  assign T124 = T125 ? io_in_3_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign T125 = T67[1'h0];
  assign T126 = T67[1'h1];
  assign T127 = T132 ? T130 : T128;
  assign T128 = T129 ? io_in_5_bits_manager_xact_id : io_in_4_bits_manager_xact_id;
  assign T129 = T67[1'h0];
  assign T130 = T131 ? io_in_7_bits_manager_xact_id : io_in_6_bits_manager_xact_id;
  assign T131 = T67[1'h0];
  assign T132 = T67[1'h1];
  assign T133 = T67[2'h2];
  assign io_out_bits_client_xact_id = T134;
  assign T134 = T147 ? T141 : T135;
  assign T135 = T140 ? T138 : T136;
  assign T136 = T137 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T137 = T67[1'h0];
  assign T138 = T139 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T139 = T67[1'h0];
  assign T140 = T67[1'h1];
  assign T141 = T146 ? T144 : T142;
  assign T142 = T143 ? io_in_5_bits_client_xact_id : io_in_4_bits_client_xact_id;
  assign T143 = T67[1'h0];
  assign T144 = T145 ? io_in_7_bits_client_xact_id : io_in_6_bits_client_xact_id;
  assign T145 = T67[1'h0];
  assign T146 = T67[1'h1];
  assign T147 = T67[2'h2];
  assign io_out_bits_addr_beat = T148;
  assign T148 = T161 ? T155 : T149;
  assign T149 = T154 ? T152 : T150;
  assign T150 = T151 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T151 = T67[1'h0];
  assign T152 = T153 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T153 = T67[1'h0];
  assign T154 = T67[1'h1];
  assign T155 = T160 ? T158 : T156;
  assign T156 = T157 ? io_in_5_bits_addr_beat : io_in_4_bits_addr_beat;
  assign T157 = T67[1'h0];
  assign T158 = T159 ? io_in_7_bits_addr_beat : io_in_6_bits_addr_beat;
  assign T159 = T67[1'h0];
  assign T160 = T67[1'h1];
  assign T161 = T67[2'h2];
  assign io_out_valid = T162;
  assign T162 = T175 ? T169 : T163;
  assign T163 = T168 ? T166 : T164;
  assign T164 = T165 ? io_in_1_valid : io_in_0_valid;
  assign T165 = T67[1'h0];
  assign T166 = T167 ? io_in_3_valid : io_in_2_valid;
  assign T167 = T67[1'h0];
  assign T168 = T67[1'h1];
  assign T169 = T174 ? T172 : T170;
  assign T170 = T171 ? io_in_5_valid : io_in_4_valid;
  assign T171 = T67[1'h0];
  assign T172 = T173 ? io_in_7_valid : io_in_6_valid;
  assign T173 = T67[1'h0];
  assign T174 = T67[1'h1];
  assign T175 = T67[2'h2];
  assign io_in_0_ready = T176;
  assign T176 = T177 & io_out_ready;
  assign T177 = locked ? T204 : T178;
  assign T178 = T203 | T179;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T183 | T181;
  assign T181 = io_in_7_valid & T182;
  assign T182 = last_grant < 3'h7;
  assign T183 = T186 | T184;
  assign T184 = io_in_6_valid & T185;
  assign T185 = last_grant < 3'h6;
  assign T186 = T189 | T187;
  assign T187 = io_in_5_valid & T188;
  assign T188 = last_grant < 3'h5;
  assign T189 = T192 | T190;
  assign T190 = io_in_4_valid & T191;
  assign T191 = last_grant < 3'h4;
  assign T192 = T195 | T193;
  assign T193 = io_in_3_valid & T194;
  assign T194 = last_grant < 3'h3;
  assign T195 = T198 | T196;
  assign T196 = io_in_2_valid & T197;
  assign T197 = last_grant < 3'h2;
  assign T198 = T201 | T199;
  assign T199 = io_in_1_valid & T200;
  assign T200 = last_grant < 3'h1;
  assign T201 = io_in_0_valid & T202;
  assign T202 = last_grant < 3'h0;
  assign T203 = last_grant < 3'h0;
  assign T204 = lockIdx == 3'h0;
  assign io_in_1_ready = T205;
  assign T205 = T206 & io_out_ready;
  assign T206 = locked ? T220 : T207;
  assign T207 = T217 | T208;
  assign T208 = T209 ^ 1'h1;
  assign T209 = T210 | io_in_0_valid;
  assign T210 = T211 | T181;
  assign T211 = T212 | T184;
  assign T212 = T213 | T187;
  assign T213 = T214 | T190;
  assign T214 = T215 | T193;
  assign T215 = T216 | T196;
  assign T216 = T201 | T199;
  assign T217 = T219 & T218;
  assign T218 = last_grant < 3'h1;
  assign T219 = T201 ^ 1'h1;
  assign T220 = lockIdx == 3'h1;
  assign io_in_2_ready = T221;
  assign T221 = T222 & io_out_ready;
  assign T222 = locked ? T238 : T223;
  assign T223 = T234 | T224;
  assign T224 = T225 ^ 1'h1;
  assign T225 = T226 | io_in_1_valid;
  assign T226 = T227 | io_in_0_valid;
  assign T227 = T228 | T181;
  assign T228 = T229 | T184;
  assign T229 = T230 | T187;
  assign T230 = T231 | T190;
  assign T231 = T232 | T193;
  assign T232 = T233 | T196;
  assign T233 = T201 | T199;
  assign T234 = T236 & T235;
  assign T235 = last_grant < 3'h2;
  assign T236 = T237 ^ 1'h1;
  assign T237 = T201 | T199;
  assign T238 = lockIdx == 3'h2;
  assign io_in_3_ready = T239;
  assign T239 = T240 & io_out_ready;
  assign T240 = locked ? T258 : T241;
  assign T241 = T253 | T242;
  assign T242 = T243 ^ 1'h1;
  assign T243 = T244 | io_in_2_valid;
  assign T244 = T245 | io_in_1_valid;
  assign T245 = T246 | io_in_0_valid;
  assign T246 = T247 | T181;
  assign T247 = T248 | T184;
  assign T248 = T249 | T187;
  assign T249 = T250 | T190;
  assign T250 = T251 | T193;
  assign T251 = T252 | T196;
  assign T252 = T201 | T199;
  assign T253 = T255 & T254;
  assign T254 = last_grant < 3'h3;
  assign T255 = T256 ^ 1'h1;
  assign T256 = T257 | T196;
  assign T257 = T201 | T199;
  assign T258 = lockIdx == 3'h3;
  assign io_in_4_ready = T259;
  assign T259 = T260 & io_out_ready;
  assign T260 = locked ? T280 : T261;
  assign T261 = T274 | T262;
  assign T262 = T263 ^ 1'h1;
  assign T263 = T264 | io_in_3_valid;
  assign T264 = T265 | io_in_2_valid;
  assign T265 = T266 | io_in_1_valid;
  assign T266 = T267 | io_in_0_valid;
  assign T267 = T268 | T181;
  assign T268 = T269 | T184;
  assign T269 = T270 | T187;
  assign T270 = T271 | T190;
  assign T271 = T272 | T193;
  assign T272 = T273 | T196;
  assign T273 = T201 | T199;
  assign T274 = T276 & T275;
  assign T275 = last_grant < 3'h4;
  assign T276 = T277 ^ 1'h1;
  assign T277 = T278 | T193;
  assign T278 = T279 | T196;
  assign T279 = T201 | T199;
  assign T280 = lockIdx == 3'h4;
  assign io_in_5_ready = T281;
  assign T281 = T282 & io_out_ready;
  assign T282 = locked ? T304 : T283;
  assign T283 = T297 | T284;
  assign T284 = T285 ^ 1'h1;
  assign T285 = T286 | io_in_4_valid;
  assign T286 = T287 | io_in_3_valid;
  assign T287 = T288 | io_in_2_valid;
  assign T288 = T289 | io_in_1_valid;
  assign T289 = T290 | io_in_0_valid;
  assign T290 = T291 | T181;
  assign T291 = T292 | T184;
  assign T292 = T293 | T187;
  assign T293 = T294 | T190;
  assign T294 = T295 | T193;
  assign T295 = T296 | T196;
  assign T296 = T201 | T199;
  assign T297 = T299 & T298;
  assign T298 = last_grant < 3'h5;
  assign T299 = T300 ^ 1'h1;
  assign T300 = T301 | T190;
  assign T301 = T302 | T193;
  assign T302 = T303 | T196;
  assign T303 = T201 | T199;
  assign T304 = lockIdx == 3'h5;
  assign io_in_6_ready = T305;
  assign T305 = T306 & io_out_ready;
  assign T306 = locked ? T330 : T307;
  assign T307 = T322 | T308;
  assign T308 = T309 ^ 1'h1;
  assign T309 = T310 | io_in_5_valid;
  assign T310 = T311 | io_in_4_valid;
  assign T311 = T312 | io_in_3_valid;
  assign T312 = T313 | io_in_2_valid;
  assign T313 = T314 | io_in_1_valid;
  assign T314 = T315 | io_in_0_valid;
  assign T315 = T316 | T181;
  assign T316 = T317 | T184;
  assign T317 = T318 | T187;
  assign T318 = T319 | T190;
  assign T319 = T320 | T193;
  assign T320 = T321 | T196;
  assign T321 = T201 | T199;
  assign T322 = T324 & T323;
  assign T323 = last_grant < 3'h6;
  assign T324 = T325 ^ 1'h1;
  assign T325 = T326 | T187;
  assign T326 = T327 | T190;
  assign T327 = T328 | T193;
  assign T328 = T329 | T196;
  assign T329 = T201 | T199;
  assign T330 = lockIdx == 3'h6;
  assign io_in_7_ready = T331;
  assign T331 = T332 & io_out_ready;
  assign T332 = locked ? T358 : T333;
  assign T333 = T349 | T334;
  assign T334 = T335 ^ 1'h1;
  assign T335 = T336 | io_in_6_valid;
  assign T336 = T337 | io_in_5_valid;
  assign T337 = T338 | io_in_4_valid;
  assign T338 = T339 | io_in_3_valid;
  assign T339 = T340 | io_in_2_valid;
  assign T340 = T341 | io_in_1_valid;
  assign T341 = T342 | io_in_0_valid;
  assign T342 = T343 | T181;
  assign T343 = T344 | T184;
  assign T344 = T345 | T187;
  assign T345 = T346 | T190;
  assign T346 = T347 | T193;
  assign T347 = T348 | T196;
  assign T348 = T201 | T199;
  assign T349 = T351 & T350;
  assign T350 = last_grant < 3'h7;
  assign T351 = T352 ^ 1'h1;
  assign T352 = T353 | T184;
  assign T353 = T354 | T187;
  assign T354 = T355 | T190;
  assign T355 = T356 | T193;
  assign T356 = T357 | T196;
  assign T357 = T201 | T199;
  assign T358 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T45) begin
      lockIdx <= T31;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T61) begin
      locked <= 1'h0;
    end else if(T47) begin
      locked <= T56;
    end
    if(reset) begin
      R59 <= 2'h0;
    end else if(T47) begin
      R59 <= T58;
    end
  end
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [25:0] io_in_7_bits_addr_block,
    input [1:0] io_in_7_bits_p_type,
    input [1:0] io_in_7_bits_client_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [25:0] io_in_6_bits_addr_block,
    input [1:0] io_in_6_bits_p_type,
    input [1:0] io_in_6_bits_client_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [25:0] io_in_5_bits_addr_block,
    input [1:0] io_in_5_bits_p_type,
    input [1:0] io_in_5_bits_client_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [1:0] io_in_4_bits_p_type,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [1:0] io_in_3_bits_p_type,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_p_type,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_p_type,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_p_type,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_p_type,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T272;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T273;
  reg  locked;
  wire T274;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[25:0] T61;
  wire[25:0] T62;
  wire[25:0] T63;
  wire T64;
  wire[25:0] T65;
  wire T66;
  wire T67;
  wire[25:0] T68;
  wire[25:0] T69;
  wire T70;
  wire[25:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T272 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T273 = reset ? 3'h7 : lockIdx;
  assign T274 = reset ? 1'h0 : T30;
  assign T30 = T31 ? 1'h0 : locked;
  assign T31 = io_out_valid & io_out_ready;
  assign io_out_bits_client_id = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T35 = T36[1'h0];
  assign T36 = chosen;
  assign T37 = T38 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T38 = T36[1'h0];
  assign T39 = T36[1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_client_id : io_in_4_bits_client_id;
  assign T42 = T36[1'h0];
  assign T43 = T44 ? io_in_7_bits_client_id : io_in_6_bits_client_id;
  assign T44 = T36[1'h0];
  assign T45 = T36[1'h1];
  assign T46 = T36[2'h2];
  assign io_out_bits_p_type = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign T50 = T36[1'h0];
  assign T51 = T52 ? io_in_3_bits_p_type : io_in_2_bits_p_type;
  assign T52 = T36[1'h0];
  assign T53 = T36[1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_p_type : io_in_4_bits_p_type;
  assign T56 = T36[1'h0];
  assign T57 = T58 ? io_in_7_bits_p_type : io_in_6_bits_p_type;
  assign T58 = T36[1'h0];
  assign T59 = T36[1'h1];
  assign T60 = T36[2'h2];
  assign io_out_bits_addr_block = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T64 = T36[1'h0];
  assign T65 = T66 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T66 = T36[1'h0];
  assign T67 = T36[1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_addr_block : io_in_4_bits_addr_block;
  assign T70 = T36[1'h0];
  assign T71 = T72 ? io_in_7_bits_addr_block : io_in_6_bits_addr_block;
  assign T72 = T36[1'h0];
  assign T73 = T36[1'h1];
  assign T74 = T36[2'h2];
  assign io_out_valid = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_valid : io_in_0_valid;
  assign T78 = T36[1'h0];
  assign T79 = T80 ? io_in_3_valid : io_in_2_valid;
  assign T80 = T36[1'h0];
  assign T81 = T36[1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_valid : io_in_4_valid;
  assign T84 = T36[1'h0];
  assign T85 = T86 ? io_in_7_valid : io_in_6_valid;
  assign T86 = T36[1'h0];
  assign T87 = T36[1'h1];
  assign T88 = T36[2'h2];
  assign io_in_0_ready = T89;
  assign T89 = T90 & io_out_ready;
  assign T90 = locked ? T117 : T91;
  assign T91 = T116 | T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T96 | T94;
  assign T94 = io_in_7_valid & T95;
  assign T95 = last_grant < 3'h7;
  assign T96 = T99 | T97;
  assign T97 = io_in_6_valid & T98;
  assign T98 = last_grant < 3'h6;
  assign T99 = T102 | T100;
  assign T100 = io_in_5_valid & T101;
  assign T101 = last_grant < 3'h5;
  assign T102 = T105 | T103;
  assign T103 = io_in_4_valid & T104;
  assign T104 = last_grant < 3'h4;
  assign T105 = T108 | T106;
  assign T106 = io_in_3_valid & T107;
  assign T107 = last_grant < 3'h3;
  assign T108 = T111 | T109;
  assign T109 = io_in_2_valid & T110;
  assign T110 = last_grant < 3'h2;
  assign T111 = T114 | T112;
  assign T112 = io_in_1_valid & T113;
  assign T113 = last_grant < 3'h1;
  assign T114 = io_in_0_valid & T115;
  assign T115 = last_grant < 3'h0;
  assign T116 = last_grant < 3'h0;
  assign T117 = lockIdx == 3'h0;
  assign io_in_1_ready = T118;
  assign T118 = T119 & io_out_ready;
  assign T119 = locked ? T133 : T120;
  assign T120 = T130 | T121;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T123 | io_in_0_valid;
  assign T123 = T124 | T94;
  assign T124 = T125 | T97;
  assign T125 = T126 | T100;
  assign T126 = T127 | T103;
  assign T127 = T128 | T106;
  assign T128 = T129 | T109;
  assign T129 = T114 | T112;
  assign T130 = T132 & T131;
  assign T131 = last_grant < 3'h1;
  assign T132 = T114 ^ 1'h1;
  assign T133 = lockIdx == 3'h1;
  assign io_in_2_ready = T134;
  assign T134 = T135 & io_out_ready;
  assign T135 = locked ? T151 : T136;
  assign T136 = T147 | T137;
  assign T137 = T138 ^ 1'h1;
  assign T138 = T139 | io_in_1_valid;
  assign T139 = T140 | io_in_0_valid;
  assign T140 = T141 | T94;
  assign T141 = T142 | T97;
  assign T142 = T143 | T100;
  assign T143 = T144 | T103;
  assign T144 = T145 | T106;
  assign T145 = T146 | T109;
  assign T146 = T114 | T112;
  assign T147 = T149 & T148;
  assign T148 = last_grant < 3'h2;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T114 | T112;
  assign T151 = lockIdx == 3'h2;
  assign io_in_3_ready = T152;
  assign T152 = T153 & io_out_ready;
  assign T153 = locked ? T171 : T154;
  assign T154 = T166 | T155;
  assign T155 = T156 ^ 1'h1;
  assign T156 = T157 | io_in_2_valid;
  assign T157 = T158 | io_in_1_valid;
  assign T158 = T159 | io_in_0_valid;
  assign T159 = T160 | T94;
  assign T160 = T161 | T97;
  assign T161 = T162 | T100;
  assign T162 = T163 | T103;
  assign T163 = T164 | T106;
  assign T164 = T165 | T109;
  assign T165 = T114 | T112;
  assign T166 = T168 & T167;
  assign T167 = last_grant < 3'h3;
  assign T168 = T169 ^ 1'h1;
  assign T169 = T170 | T109;
  assign T170 = T114 | T112;
  assign T171 = lockIdx == 3'h3;
  assign io_in_4_ready = T172;
  assign T172 = T173 & io_out_ready;
  assign T173 = locked ? T193 : T174;
  assign T174 = T187 | T175;
  assign T175 = T176 ^ 1'h1;
  assign T176 = T177 | io_in_3_valid;
  assign T177 = T178 | io_in_2_valid;
  assign T178 = T179 | io_in_1_valid;
  assign T179 = T180 | io_in_0_valid;
  assign T180 = T181 | T94;
  assign T181 = T182 | T97;
  assign T182 = T183 | T100;
  assign T183 = T184 | T103;
  assign T184 = T185 | T106;
  assign T185 = T186 | T109;
  assign T186 = T114 | T112;
  assign T187 = T189 & T188;
  assign T188 = last_grant < 3'h4;
  assign T189 = T190 ^ 1'h1;
  assign T190 = T191 | T106;
  assign T191 = T192 | T109;
  assign T192 = T114 | T112;
  assign T193 = lockIdx == 3'h4;
  assign io_in_5_ready = T194;
  assign T194 = T195 & io_out_ready;
  assign T195 = locked ? T217 : T196;
  assign T196 = T210 | T197;
  assign T197 = T198 ^ 1'h1;
  assign T198 = T199 | io_in_4_valid;
  assign T199 = T200 | io_in_3_valid;
  assign T200 = T201 | io_in_2_valid;
  assign T201 = T202 | io_in_1_valid;
  assign T202 = T203 | io_in_0_valid;
  assign T203 = T204 | T94;
  assign T204 = T205 | T97;
  assign T205 = T206 | T100;
  assign T206 = T207 | T103;
  assign T207 = T208 | T106;
  assign T208 = T209 | T109;
  assign T209 = T114 | T112;
  assign T210 = T212 & T211;
  assign T211 = last_grant < 3'h5;
  assign T212 = T213 ^ 1'h1;
  assign T213 = T214 | T103;
  assign T214 = T215 | T106;
  assign T215 = T216 | T109;
  assign T216 = T114 | T112;
  assign T217 = lockIdx == 3'h5;
  assign io_in_6_ready = T218;
  assign T218 = T219 & io_out_ready;
  assign T219 = locked ? T243 : T220;
  assign T220 = T235 | T221;
  assign T221 = T222 ^ 1'h1;
  assign T222 = T223 | io_in_5_valid;
  assign T223 = T224 | io_in_4_valid;
  assign T224 = T225 | io_in_3_valid;
  assign T225 = T226 | io_in_2_valid;
  assign T226 = T227 | io_in_1_valid;
  assign T227 = T228 | io_in_0_valid;
  assign T228 = T229 | T94;
  assign T229 = T230 | T97;
  assign T230 = T231 | T100;
  assign T231 = T232 | T103;
  assign T232 = T233 | T106;
  assign T233 = T234 | T109;
  assign T234 = T114 | T112;
  assign T235 = T237 & T236;
  assign T236 = last_grant < 3'h6;
  assign T237 = T238 ^ 1'h1;
  assign T238 = T239 | T100;
  assign T239 = T240 | T103;
  assign T240 = T241 | T106;
  assign T241 = T242 | T109;
  assign T242 = T114 | T112;
  assign T243 = lockIdx == 3'h6;
  assign io_in_7_ready = T244;
  assign T244 = T245 & io_out_ready;
  assign T245 = locked ? T271 : T246;
  assign T246 = T262 | T247;
  assign T247 = T248 ^ 1'h1;
  assign T248 = T249 | io_in_6_valid;
  assign T249 = T250 | io_in_5_valid;
  assign T250 = T251 | io_in_4_valid;
  assign T251 = T252 | io_in_3_valid;
  assign T252 = T253 | io_in_2_valid;
  assign T253 = T254 | io_in_1_valid;
  assign T254 = T255 | io_in_0_valid;
  assign T255 = T256 | T94;
  assign T256 = T257 | T97;
  assign T257 = T258 | T100;
  assign T258 = T259 | T103;
  assign T259 = T260 | T106;
  assign T260 = T261 | T109;
  assign T261 = T114 | T112;
  assign T262 = T264 & T263;
  assign T263 = last_grant < 3'h7;
  assign T264 = T265 ^ 1'h1;
  assign T265 = T266 | T97;
  assign T266 = T267 | T100;
  assign T267 = T268 | T103;
  assign T268 = T269 | T106;
  assign T269 = T270 | T109;
  assign T270 = T114 | T112;
  assign T271 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T31) begin
      locked <= 1'h0;
    end
  end
endmodule

module LockingRRArbiter_10(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [25:0] io_in_7_bits_addr_block,
    input [3:0] io_in_7_bits_client_xact_id,
    input [1:0] io_in_7_bits_addr_beat,
    input  io_in_7_bits_is_builtin_type,
    input [2:0] io_in_7_bits_a_type,
    input [16:0] io_in_7_bits_union,
    input [3:0] io_in_7_bits_data,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [25:0] io_in_6_bits_addr_block,
    input [3:0] io_in_6_bits_client_xact_id,
    input [1:0] io_in_6_bits_addr_beat,
    input  io_in_6_bits_is_builtin_type,
    input [2:0] io_in_6_bits_a_type,
    input [16:0] io_in_6_bits_union,
    input [3:0] io_in_6_bits_data,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [25:0] io_in_5_bits_addr_block,
    input [3:0] io_in_5_bits_client_xact_id,
    input [1:0] io_in_5_bits_addr_beat,
    input  io_in_5_bits_is_builtin_type,
    input [2:0] io_in_5_bits_a_type,
    input [16:0] io_in_5_bits_union,
    input [3:0] io_in_5_bits_data,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [3:0] io_in_4_bits_client_xact_id,
    input [1:0] io_in_4_bits_addr_beat,
    input  io_in_4_bits_is_builtin_type,
    input [2:0] io_in_4_bits_a_type,
    input [16:0] io_in_4_bits_union,
    input [3:0] io_in_4_bits_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [3:0] io_in_3_bits_client_xact_id,
    input [1:0] io_in_3_bits_addr_beat,
    input  io_in_3_bits_is_builtin_type,
    input [2:0] io_in_3_bits_a_type,
    input [16:0] io_in_3_bits_union,
    input [3:0] io_in_3_bits_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [3:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [3:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [3:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [3:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [3:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [3:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[3:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[3:0] io_out_bits_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T356;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T357;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  locked;
  wire T358;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  reg [1:0] R56;
  wire[1:0] T359;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire T63;
  wire[2:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire[3:0] T68;
  wire[3:0] T69;
  wire T70;
  wire[3:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[16:0] T75;
  wire[16:0] T76;
  wire[16:0] T77;
  wire T78;
  wire[16:0] T79;
  wire T80;
  wire T81;
  wire[16:0] T82;
  wire[16:0] T83;
  wire T84;
  wire[16:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire[2:0] T90;
  wire[2:0] T91;
  wire T92;
  wire[2:0] T93;
  wire T94;
  wire T95;
  wire[2:0] T96;
  wire[2:0] T97;
  wire T98;
  wire[2:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire[1:0] T121;
  wire T122;
  wire T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire T126;
  wire[1:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[3:0] T131;
  wire[3:0] T132;
  wire[3:0] T133;
  wire T134;
  wire[3:0] T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[25:0] T145;
  wire[25:0] T146;
  wire[25:0] T147;
  wire T148;
  wire[25:0] T149;
  wire T150;
  wire T151;
  wire[25:0] T152;
  wire[25:0] T153;
  wire T154;
  wire[25:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R56 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T356 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T357 = reset ? 3'h7 : T30;
  assign T30 = T45 ? T31 : lockIdx;
  assign T31 = T44 ? 3'h0 : T32;
  assign T32 = T43 ? 3'h1 : T33;
  assign T33 = T42 ? 3'h2 : T34;
  assign T34 = T41 ? 3'h3 : T35;
  assign T35 = T40 ? 3'h4 : T36;
  assign T36 = T39 ? 3'h5 : T37;
  assign T37 = T38 ? 3'h6 : 3'h7;
  assign T38 = io_in_6_ready & io_in_6_valid;
  assign T39 = io_in_5_ready & io_in_5_valid;
  assign T40 = io_in_4_ready & io_in_4_valid;
  assign T41 = io_in_3_ready & io_in_3_valid;
  assign T42 = io_in_2_ready & io_in_2_valid;
  assign T43 = io_in_1_ready & io_in_1_valid;
  assign T44 = io_in_0_ready & io_in_0_valid;
  assign T45 = T47 & T46;
  assign T46 = locked ^ 1'h1;
  assign T47 = T50 & T48;
  assign T48 = io_out_bits_is_builtin_type & T49;
  assign T49 = 3'h3 == io_out_bits_a_type;
  assign T50 = io_out_valid & io_out_ready;
  assign T358 = reset ? 1'h0 : T51;
  assign T51 = T58 ? 1'h0 : T52;
  assign T52 = T47 ? T53 : locked;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T55 == 2'h0;
  assign T55 = R56 + 2'h1;
  assign T359 = reset ? 2'h0 : T57;
  assign T57 = T47 ? T55 : R56;
  assign T58 = T50 & T59;
  assign T59 = T48 ^ 1'h1;
  assign io_out_bits_data = T60;
  assign T60 = T74 ? T68 : T61;
  assign T61 = T67 ? T65 : T62;
  assign T62 = T63 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T63 = T64[1'h0];
  assign T64 = chosen;
  assign T65 = T66 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T66 = T64[1'h0];
  assign T67 = T64[1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_data : io_in_4_bits_data;
  assign T70 = T64[1'h0];
  assign T71 = T72 ? io_in_7_bits_data : io_in_6_bits_data;
  assign T72 = T64[1'h0];
  assign T73 = T64[1'h1];
  assign T74 = T64[2'h2];
  assign io_out_bits_union = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T78 = T64[1'h0];
  assign T79 = T80 ? io_in_3_bits_union : io_in_2_bits_union;
  assign T80 = T64[1'h0];
  assign T81 = T64[1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_bits_union : io_in_4_bits_union;
  assign T84 = T64[1'h0];
  assign T85 = T86 ? io_in_7_bits_union : io_in_6_bits_union;
  assign T86 = T64[1'h0];
  assign T87 = T64[1'h1];
  assign T88 = T64[2'h2];
  assign io_out_bits_a_type = T89;
  assign T89 = T102 ? T96 : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T92 = T64[1'h0];
  assign T93 = T94 ? io_in_3_bits_a_type : io_in_2_bits_a_type;
  assign T94 = T64[1'h0];
  assign T95 = T64[1'h1];
  assign T96 = T101 ? T99 : T97;
  assign T97 = T98 ? io_in_5_bits_a_type : io_in_4_bits_a_type;
  assign T98 = T64[1'h0];
  assign T99 = T100 ? io_in_7_bits_a_type : io_in_6_bits_a_type;
  assign T100 = T64[1'h0];
  assign T101 = T64[1'h1];
  assign T102 = T64[2'h2];
  assign io_out_bits_is_builtin_type = T103;
  assign T103 = T116 ? T110 : T104;
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T106 = T64[1'h0];
  assign T107 = T108 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T108 = T64[1'h0];
  assign T109 = T64[1'h1];
  assign T110 = T115 ? T113 : T111;
  assign T111 = T112 ? io_in_5_bits_is_builtin_type : io_in_4_bits_is_builtin_type;
  assign T112 = T64[1'h0];
  assign T113 = T114 ? io_in_7_bits_is_builtin_type : io_in_6_bits_is_builtin_type;
  assign T114 = T64[1'h0];
  assign T115 = T64[1'h1];
  assign T116 = T64[2'h2];
  assign io_out_bits_addr_beat = T117;
  assign T117 = T130 ? T124 : T118;
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T120 = T64[1'h0];
  assign T121 = T122 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T122 = T64[1'h0];
  assign T123 = T64[1'h1];
  assign T124 = T129 ? T127 : T125;
  assign T125 = T126 ? io_in_5_bits_addr_beat : io_in_4_bits_addr_beat;
  assign T126 = T64[1'h0];
  assign T127 = T128 ? io_in_7_bits_addr_beat : io_in_6_bits_addr_beat;
  assign T128 = T64[1'h0];
  assign T129 = T64[1'h1];
  assign T130 = T64[2'h2];
  assign io_out_bits_client_xact_id = T131;
  assign T131 = T144 ? T138 : T132;
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T134 = T64[1'h0];
  assign T135 = T136 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T136 = T64[1'h0];
  assign T137 = T64[1'h1];
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140 ? io_in_5_bits_client_xact_id : io_in_4_bits_client_xact_id;
  assign T140 = T64[1'h0];
  assign T141 = T142 ? io_in_7_bits_client_xact_id : io_in_6_bits_client_xact_id;
  assign T142 = T64[1'h0];
  assign T143 = T64[1'h1];
  assign T144 = T64[2'h2];
  assign io_out_bits_addr_block = T145;
  assign T145 = T158 ? T152 : T146;
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T148 = T64[1'h0];
  assign T149 = T150 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T150 = T64[1'h0];
  assign T151 = T64[1'h1];
  assign T152 = T157 ? T155 : T153;
  assign T153 = T154 ? io_in_5_bits_addr_block : io_in_4_bits_addr_block;
  assign T154 = T64[1'h0];
  assign T155 = T156 ? io_in_7_bits_addr_block : io_in_6_bits_addr_block;
  assign T156 = T64[1'h0];
  assign T157 = T64[1'h1];
  assign T158 = T64[2'h2];
  assign io_out_valid = T159;
  assign T159 = T172 ? T166 : T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162 ? io_in_1_valid : io_in_0_valid;
  assign T162 = T64[1'h0];
  assign T163 = T164 ? io_in_3_valid : io_in_2_valid;
  assign T164 = T64[1'h0];
  assign T165 = T64[1'h1];
  assign T166 = T171 ? T169 : T167;
  assign T167 = T168 ? io_in_5_valid : io_in_4_valid;
  assign T168 = T64[1'h0];
  assign T169 = T170 ? io_in_7_valid : io_in_6_valid;
  assign T170 = T64[1'h0];
  assign T171 = T64[1'h1];
  assign T172 = T64[2'h2];
  assign io_in_0_ready = T173;
  assign T173 = T174 & io_out_ready;
  assign T174 = locked ? T201 : T175;
  assign T175 = T200 | T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T180 | T178;
  assign T178 = io_in_7_valid & T179;
  assign T179 = last_grant < 3'h7;
  assign T180 = T183 | T181;
  assign T181 = io_in_6_valid & T182;
  assign T182 = last_grant < 3'h6;
  assign T183 = T186 | T184;
  assign T184 = io_in_5_valid & T185;
  assign T185 = last_grant < 3'h5;
  assign T186 = T189 | T187;
  assign T187 = io_in_4_valid & T188;
  assign T188 = last_grant < 3'h4;
  assign T189 = T192 | T190;
  assign T190 = io_in_3_valid & T191;
  assign T191 = last_grant < 3'h3;
  assign T192 = T195 | T193;
  assign T193 = io_in_2_valid & T194;
  assign T194 = last_grant < 3'h2;
  assign T195 = T198 | T196;
  assign T196 = io_in_1_valid & T197;
  assign T197 = last_grant < 3'h1;
  assign T198 = io_in_0_valid & T199;
  assign T199 = last_grant < 3'h0;
  assign T200 = last_grant < 3'h0;
  assign T201 = lockIdx == 3'h0;
  assign io_in_1_ready = T202;
  assign T202 = T203 & io_out_ready;
  assign T203 = locked ? T217 : T204;
  assign T204 = T214 | T205;
  assign T205 = T206 ^ 1'h1;
  assign T206 = T207 | io_in_0_valid;
  assign T207 = T208 | T178;
  assign T208 = T209 | T181;
  assign T209 = T210 | T184;
  assign T210 = T211 | T187;
  assign T211 = T212 | T190;
  assign T212 = T213 | T193;
  assign T213 = T198 | T196;
  assign T214 = T216 & T215;
  assign T215 = last_grant < 3'h1;
  assign T216 = T198 ^ 1'h1;
  assign T217 = lockIdx == 3'h1;
  assign io_in_2_ready = T218;
  assign T218 = T219 & io_out_ready;
  assign T219 = locked ? T235 : T220;
  assign T220 = T231 | T221;
  assign T221 = T222 ^ 1'h1;
  assign T222 = T223 | io_in_1_valid;
  assign T223 = T224 | io_in_0_valid;
  assign T224 = T225 | T178;
  assign T225 = T226 | T181;
  assign T226 = T227 | T184;
  assign T227 = T228 | T187;
  assign T228 = T229 | T190;
  assign T229 = T230 | T193;
  assign T230 = T198 | T196;
  assign T231 = T233 & T232;
  assign T232 = last_grant < 3'h2;
  assign T233 = T234 ^ 1'h1;
  assign T234 = T198 | T196;
  assign T235 = lockIdx == 3'h2;
  assign io_in_3_ready = T236;
  assign T236 = T237 & io_out_ready;
  assign T237 = locked ? T255 : T238;
  assign T238 = T250 | T239;
  assign T239 = T240 ^ 1'h1;
  assign T240 = T241 | io_in_2_valid;
  assign T241 = T242 | io_in_1_valid;
  assign T242 = T243 | io_in_0_valid;
  assign T243 = T244 | T178;
  assign T244 = T245 | T181;
  assign T245 = T246 | T184;
  assign T246 = T247 | T187;
  assign T247 = T248 | T190;
  assign T248 = T249 | T193;
  assign T249 = T198 | T196;
  assign T250 = T252 & T251;
  assign T251 = last_grant < 3'h3;
  assign T252 = T253 ^ 1'h1;
  assign T253 = T254 | T193;
  assign T254 = T198 | T196;
  assign T255 = lockIdx == 3'h3;
  assign io_in_4_ready = T256;
  assign T256 = T257 & io_out_ready;
  assign T257 = locked ? T277 : T258;
  assign T258 = T271 | T259;
  assign T259 = T260 ^ 1'h1;
  assign T260 = T261 | io_in_3_valid;
  assign T261 = T262 | io_in_2_valid;
  assign T262 = T263 | io_in_1_valid;
  assign T263 = T264 | io_in_0_valid;
  assign T264 = T265 | T178;
  assign T265 = T266 | T181;
  assign T266 = T267 | T184;
  assign T267 = T268 | T187;
  assign T268 = T269 | T190;
  assign T269 = T270 | T193;
  assign T270 = T198 | T196;
  assign T271 = T273 & T272;
  assign T272 = last_grant < 3'h4;
  assign T273 = T274 ^ 1'h1;
  assign T274 = T275 | T190;
  assign T275 = T276 | T193;
  assign T276 = T198 | T196;
  assign T277 = lockIdx == 3'h4;
  assign io_in_5_ready = T278;
  assign T278 = T279 & io_out_ready;
  assign T279 = locked ? T301 : T280;
  assign T280 = T294 | T281;
  assign T281 = T282 ^ 1'h1;
  assign T282 = T283 | io_in_4_valid;
  assign T283 = T284 | io_in_3_valid;
  assign T284 = T285 | io_in_2_valid;
  assign T285 = T286 | io_in_1_valid;
  assign T286 = T287 | io_in_0_valid;
  assign T287 = T288 | T178;
  assign T288 = T289 | T181;
  assign T289 = T290 | T184;
  assign T290 = T291 | T187;
  assign T291 = T292 | T190;
  assign T292 = T293 | T193;
  assign T293 = T198 | T196;
  assign T294 = T296 & T295;
  assign T295 = last_grant < 3'h5;
  assign T296 = T297 ^ 1'h1;
  assign T297 = T298 | T187;
  assign T298 = T299 | T190;
  assign T299 = T300 | T193;
  assign T300 = T198 | T196;
  assign T301 = lockIdx == 3'h5;
  assign io_in_6_ready = T302;
  assign T302 = T303 & io_out_ready;
  assign T303 = locked ? T327 : T304;
  assign T304 = T319 | T305;
  assign T305 = T306 ^ 1'h1;
  assign T306 = T307 | io_in_5_valid;
  assign T307 = T308 | io_in_4_valid;
  assign T308 = T309 | io_in_3_valid;
  assign T309 = T310 | io_in_2_valid;
  assign T310 = T311 | io_in_1_valid;
  assign T311 = T312 | io_in_0_valid;
  assign T312 = T313 | T178;
  assign T313 = T314 | T181;
  assign T314 = T315 | T184;
  assign T315 = T316 | T187;
  assign T316 = T317 | T190;
  assign T317 = T318 | T193;
  assign T318 = T198 | T196;
  assign T319 = T321 & T320;
  assign T320 = last_grant < 3'h6;
  assign T321 = T322 ^ 1'h1;
  assign T322 = T323 | T184;
  assign T323 = T324 | T187;
  assign T324 = T325 | T190;
  assign T325 = T326 | T193;
  assign T326 = T198 | T196;
  assign T327 = lockIdx == 3'h6;
  assign io_in_7_ready = T328;
  assign T328 = T329 & io_out_ready;
  assign T329 = locked ? T355 : T330;
  assign T330 = T346 | T331;
  assign T331 = T332 ^ 1'h1;
  assign T332 = T333 | io_in_6_valid;
  assign T333 = T334 | io_in_5_valid;
  assign T334 = T335 | io_in_4_valid;
  assign T335 = T336 | io_in_3_valid;
  assign T336 = T337 | io_in_2_valid;
  assign T337 = T338 | io_in_1_valid;
  assign T338 = T339 | io_in_0_valid;
  assign T339 = T340 | T178;
  assign T340 = T341 | T181;
  assign T341 = T342 | T184;
  assign T342 = T343 | T187;
  assign T343 = T344 | T190;
  assign T344 = T345 | T193;
  assign T345 = T198 | T196;
  assign T346 = T348 & T347;
  assign T347 = last_grant < 3'h7;
  assign T348 = T349 ^ 1'h1;
  assign T349 = T350 | T181;
  assign T350 = T351 | T184;
  assign T351 = T352 | T187;
  assign T352 = T353 | T190;
  assign T353 = T354 | T193;
  assign T354 = T198 | T196;
  assign T355 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T45) begin
      lockIdx <= T31;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T58) begin
      locked <= 1'h0;
    end else if(T47) begin
      locked <= T53;
    end
    if(reset) begin
      R56 <= 2'h0;
    end else if(T47) begin
      R56 <= T55;
    end
  end
endmodule

module ClientUncachedTileLinkIOArbiter(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [25:0] io_in_7_acquire_bits_addr_block,
    input [3:0] io_in_7_acquire_bits_client_xact_id,
    input [1:0] io_in_7_acquire_bits_addr_beat,
    input  io_in_7_acquire_bits_is_builtin_type,
    input [2:0] io_in_7_acquire_bits_a_type,
    input [16:0] io_in_7_acquire_bits_union,
    input [3:0] io_in_7_acquire_bits_data,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_addr_beat,
    output[3:0] io_in_7_grant_bits_client_xact_id,
    output io_in_7_grant_bits_manager_xact_id,
    output io_in_7_grant_bits_is_builtin_type,
    output[3:0] io_in_7_grant_bits_g_type,
    output[3:0] io_in_7_grant_bits_data,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [25:0] io_in_6_acquire_bits_addr_block,
    input [3:0] io_in_6_acquire_bits_client_xact_id,
    input [1:0] io_in_6_acquire_bits_addr_beat,
    input  io_in_6_acquire_bits_is_builtin_type,
    input [2:0] io_in_6_acquire_bits_a_type,
    input [16:0] io_in_6_acquire_bits_union,
    input [3:0] io_in_6_acquire_bits_data,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_addr_beat,
    output[3:0] io_in_6_grant_bits_client_xact_id,
    output io_in_6_grant_bits_manager_xact_id,
    output io_in_6_grant_bits_is_builtin_type,
    output[3:0] io_in_6_grant_bits_g_type,
    output[3:0] io_in_6_grant_bits_data,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [25:0] io_in_5_acquire_bits_addr_block,
    input [3:0] io_in_5_acquire_bits_client_xact_id,
    input [1:0] io_in_5_acquire_bits_addr_beat,
    input  io_in_5_acquire_bits_is_builtin_type,
    input [2:0] io_in_5_acquire_bits_a_type,
    input [16:0] io_in_5_acquire_bits_union,
    input [3:0] io_in_5_acquire_bits_data,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_addr_beat,
    output[3:0] io_in_5_grant_bits_client_xact_id,
    output io_in_5_grant_bits_manager_xact_id,
    output io_in_5_grant_bits_is_builtin_type,
    output[3:0] io_in_5_grant_bits_g_type,
    output[3:0] io_in_5_grant_bits_data,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [25:0] io_in_4_acquire_bits_addr_block,
    input [3:0] io_in_4_acquire_bits_client_xact_id,
    input [1:0] io_in_4_acquire_bits_addr_beat,
    input  io_in_4_acquire_bits_is_builtin_type,
    input [2:0] io_in_4_acquire_bits_a_type,
    input [16:0] io_in_4_acquire_bits_union,
    input [3:0] io_in_4_acquire_bits_data,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_addr_beat,
    output[3:0] io_in_4_grant_bits_client_xact_id,
    output io_in_4_grant_bits_manager_xact_id,
    output io_in_4_grant_bits_is_builtin_type,
    output[3:0] io_in_4_grant_bits_g_type,
    output[3:0] io_in_4_grant_bits_data,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [25:0] io_in_3_acquire_bits_addr_block,
    input [3:0] io_in_3_acquire_bits_client_xact_id,
    input [1:0] io_in_3_acquire_bits_addr_beat,
    input  io_in_3_acquire_bits_is_builtin_type,
    input [2:0] io_in_3_acquire_bits_a_type,
    input [16:0] io_in_3_acquire_bits_union,
    input [3:0] io_in_3_acquire_bits_data,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_addr_beat,
    output[3:0] io_in_3_grant_bits_client_xact_id,
    output io_in_3_grant_bits_manager_xact_id,
    output io_in_3_grant_bits_is_builtin_type,
    output[3:0] io_in_3_grant_bits_g_type,
    output[3:0] io_in_3_grant_bits_data,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [25:0] io_in_2_acquire_bits_addr_block,
    input [3:0] io_in_2_acquire_bits_client_xact_id,
    input [1:0] io_in_2_acquire_bits_addr_beat,
    input  io_in_2_acquire_bits_is_builtin_type,
    input [2:0] io_in_2_acquire_bits_a_type,
    input [16:0] io_in_2_acquire_bits_union,
    input [3:0] io_in_2_acquire_bits_data,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_addr_beat,
    output[3:0] io_in_2_grant_bits_client_xact_id,
    output io_in_2_grant_bits_manager_xact_id,
    output io_in_2_grant_bits_is_builtin_type,
    output[3:0] io_in_2_grant_bits_g_type,
    output[3:0] io_in_2_grant_bits_data,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [25:0] io_in_1_acquire_bits_addr_block,
    input [3:0] io_in_1_acquire_bits_client_xact_id,
    input [1:0] io_in_1_acquire_bits_addr_beat,
    input  io_in_1_acquire_bits_is_builtin_type,
    input [2:0] io_in_1_acquire_bits_a_type,
    input [16:0] io_in_1_acquire_bits_union,
    input [3:0] io_in_1_acquire_bits_data,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_addr_beat,
    output[3:0] io_in_1_grant_bits_client_xact_id,
    output io_in_1_grant_bits_manager_xact_id,
    output io_in_1_grant_bits_is_builtin_type,
    output[3:0] io_in_1_grant_bits_g_type,
    output[3:0] io_in_1_grant_bits_data,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [25:0] io_in_0_acquire_bits_addr_block,
    input [3:0] io_in_0_acquire_bits_client_xact_id,
    input [1:0] io_in_0_acquire_bits_addr_beat,
    input  io_in_0_acquire_bits_is_builtin_type,
    input [2:0] io_in_0_acquire_bits_a_type,
    input [16:0] io_in_0_acquire_bits_union,
    input [3:0] io_in_0_acquire_bits_data,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_addr_beat,
    output[3:0] io_in_0_grant_bits_client_xact_id,
    output io_in_0_grant_bits_manager_xact_id,
    output io_in_0_grant_bits_is_builtin_type,
    output[3:0] io_in_0_grant_bits_g_type,
    output[3:0] io_in_0_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[3:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [3:0] io_out_grant_bits_data
);

  wire[3:0] T56;
  wire[6:0] T0;
  wire[3:0] T57;
  wire[6:0] T1;
  wire[3:0] T58;
  wire[6:0] T2;
  wire[3:0] T59;
  wire[6:0] T3;
  wire[3:0] T60;
  wire[6:0] T4;
  wire[3:0] T61;
  wire[6:0] T5;
  wire[3:0] T62;
  wire[6:0] T6;
  wire[3:0] T63;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire T37;
  wire[2:0] T38;
  wire[2:0] T39;
  wire[3:0] T64;
  wire T40;
  wire T41;
  wire[3:0] T65;
  wire T42;
  wire T43;
  wire[3:0] T66;
  wire T44;
  wire T45;
  wire[3:0] T67;
  wire T46;
  wire T47;
  wire[3:0] T68;
  wire T48;
  wire T49;
  wire[3:0] T69;
  wire T50;
  wire T51;
  wire[3:0] T70;
  wire T52;
  wire T53;
  wire[3:0] T71;
  wire T54;
  wire T55;
  wire LockingRRArbiter_io_in_7_ready;
  wire LockingRRArbiter_io_in_6_ready;
  wire LockingRRArbiter_io_in_5_ready;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[25:0] LockingRRArbiter_io_out_bits_addr_block;
  wire[3:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_addr_beat;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_union;
  wire[3:0] LockingRRArbiter_io_out_bits_data;


  assign T56 = T0[2'h3:1'h0];
  assign T0 = {io_in_0_acquire_bits_client_xact_id, 3'h0};
  assign T57 = T1[2'h3:1'h0];
  assign T1 = {io_in_1_acquire_bits_client_xact_id, 3'h1};
  assign T58 = T2[2'h3:1'h0];
  assign T2 = {io_in_2_acquire_bits_client_xact_id, 3'h2};
  assign T59 = T3[2'h3:1'h0];
  assign T3 = {io_in_3_acquire_bits_client_xact_id, 3'h3};
  assign T60 = T4[2'h3:1'h0];
  assign T4 = {io_in_4_acquire_bits_client_xact_id, 3'h4};
  assign T61 = T5[2'h3:1'h0];
  assign T5 = {io_in_5_acquire_bits_client_xact_id, 3'h5};
  assign T62 = T6[2'h3:1'h0];
  assign T6 = {io_in_6_acquire_bits_client_xact_id, 3'h6};
  assign T63 = T7[2'h3:1'h0];
  assign T7 = {io_in_7_acquire_bits_client_xact_id, 3'h7};
  assign io_out_grant_ready = T8;
  assign T8 = T37 ? io_in_7_grant_ready : T9;
  assign T9 = T34 ? io_in_6_grant_ready : T10;
  assign T10 = T31 ? io_in_5_grant_ready : T11;
  assign T11 = T28 ? io_in_4_grant_ready : T12;
  assign T12 = T25 ? io_in_3_grant_ready : T13;
  assign T13 = T22 ? io_in_2_grant_ready : T14;
  assign T14 = T19 ? io_in_1_grant_ready : T15;
  assign T15 = T16 ? io_in_0_grant_ready : 1'h0;
  assign T16 = T17 == 3'h0;
  assign T17 = T18;
  assign T18 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T19 = T20 == 3'h1;
  assign T20 = T21;
  assign T21 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T22 = T23 == 3'h2;
  assign T23 = T24;
  assign T24 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T25 = T26 == 3'h3;
  assign T26 = T27;
  assign T27 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T28 = T29 == 3'h4;
  assign T29 = T30;
  assign T30 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T31 = T32 == 3'h5;
  assign T32 = T33;
  assign T33 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T34 = T35 == 3'h6;
  assign T35 = T36;
  assign T36 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign T37 = T38 == 3'h7;
  assign T38 = T39;
  assign T39 = io_out_grant_bits_client_xact_id[2'h2:1'h0];
  assign io_out_acquire_bits_data = LockingRRArbiter_io_out_bits_data;
  assign io_out_acquire_bits_union = LockingRRArbiter_io_out_bits_union;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_io_out_bits_addr_block;
  assign io_out_acquire_valid = LockingRRArbiter_io_out_valid;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_client_xact_id = T64;
  assign T64 = {3'h0, T40};
  assign T40 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_valid = T41;
  assign T41 = T16 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_io_in_0_ready;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_client_xact_id = T65;
  assign T65 = {3'h0, T42};
  assign T42 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_valid = T43;
  assign T43 = T19 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_io_in_1_ready;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_client_xact_id = T66;
  assign T66 = {3'h0, T44};
  assign T44 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_valid = T45;
  assign T45 = T22 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = LockingRRArbiter_io_in_2_ready;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_client_xact_id = T67;
  assign T67 = {3'h0, T46};
  assign T46 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_valid = T47;
  assign T47 = T25 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = LockingRRArbiter_io_in_3_ready;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_client_xact_id = T68;
  assign T68 = {3'h0, T48};
  assign T48 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_valid = T49;
  assign T49 = T28 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = LockingRRArbiter_io_in_4_ready;
  assign io_in_5_grant_bits_data = io_out_grant_bits_data;
  assign io_in_5_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_5_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_5_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_5_grant_bits_client_xact_id = T69;
  assign T69 = {3'h0, T50};
  assign T50 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_5_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_5_grant_valid = T51;
  assign T51 = T31 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = LockingRRArbiter_io_in_5_ready;
  assign io_in_6_grant_bits_data = io_out_grant_bits_data;
  assign io_in_6_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_6_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_6_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_6_grant_bits_client_xact_id = T70;
  assign T70 = {3'h0, T52};
  assign T52 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_6_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_6_grant_valid = T53;
  assign T53 = T34 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = LockingRRArbiter_io_in_6_ready;
  assign io_in_7_grant_bits_data = io_out_grant_bits_data;
  assign io_in_7_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_7_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_7_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_7_grant_bits_client_xact_id = T71;
  assign T71 = {3'h0, T54};
  assign T54 = io_out_grant_bits_client_xact_id >> 2'h3;
  assign io_in_7_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_7_grant_valid = T55;
  assign T55 = T37 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = LockingRRArbiter_io_in_7_ready;
  LockingRRArbiter_10 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_addr_block( io_in_7_acquire_bits_addr_block ),
       .io_in_7_bits_client_xact_id( T63 ),
       .io_in_7_bits_addr_beat( io_in_7_acquire_bits_addr_beat ),
       .io_in_7_bits_is_builtin_type( io_in_7_acquire_bits_is_builtin_type ),
       .io_in_7_bits_a_type( io_in_7_acquire_bits_a_type ),
       .io_in_7_bits_union( io_in_7_acquire_bits_union ),
       .io_in_7_bits_data( io_in_7_acquire_bits_data ),
       .io_in_6_ready( LockingRRArbiter_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_addr_block( io_in_6_acquire_bits_addr_block ),
       .io_in_6_bits_client_xact_id( T62 ),
       .io_in_6_bits_addr_beat( io_in_6_acquire_bits_addr_beat ),
       .io_in_6_bits_is_builtin_type( io_in_6_acquire_bits_is_builtin_type ),
       .io_in_6_bits_a_type( io_in_6_acquire_bits_a_type ),
       .io_in_6_bits_union( io_in_6_acquire_bits_union ),
       .io_in_6_bits_data( io_in_6_acquire_bits_data ),
       .io_in_5_ready( LockingRRArbiter_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_addr_block( io_in_5_acquire_bits_addr_block ),
       .io_in_5_bits_client_xact_id( T61 ),
       .io_in_5_bits_addr_beat( io_in_5_acquire_bits_addr_beat ),
       .io_in_5_bits_is_builtin_type( io_in_5_acquire_bits_is_builtin_type ),
       .io_in_5_bits_a_type( io_in_5_acquire_bits_a_type ),
       .io_in_5_bits_union( io_in_5_acquire_bits_union ),
       .io_in_5_bits_data( io_in_5_acquire_bits_data ),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_addr_block( io_in_4_acquire_bits_addr_block ),
       .io_in_4_bits_client_xact_id( T60 ),
       .io_in_4_bits_addr_beat( io_in_4_acquire_bits_addr_beat ),
       .io_in_4_bits_is_builtin_type( io_in_4_acquire_bits_is_builtin_type ),
       .io_in_4_bits_a_type( io_in_4_acquire_bits_a_type ),
       .io_in_4_bits_union( io_in_4_acquire_bits_union ),
       .io_in_4_bits_data( io_in_4_acquire_bits_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_addr_block( io_in_3_acquire_bits_addr_block ),
       .io_in_3_bits_client_xact_id( T59 ),
       .io_in_3_bits_addr_beat( io_in_3_acquire_bits_addr_beat ),
       .io_in_3_bits_is_builtin_type( io_in_3_acquire_bits_is_builtin_type ),
       .io_in_3_bits_a_type( io_in_3_acquire_bits_a_type ),
       .io_in_3_bits_union( io_in_3_acquire_bits_union ),
       .io_in_3_bits_data( io_in_3_acquire_bits_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_addr_block( io_in_2_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( T58 ),
       .io_in_2_bits_addr_beat( io_in_2_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( io_in_2_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( io_in_2_acquire_bits_a_type ),
       .io_in_2_bits_union( io_in_2_acquire_bits_union ),
       .io_in_2_bits_data( io_in_2_acquire_bits_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_addr_block( io_in_1_acquire_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T57 ),
       .io_in_1_bits_addr_beat( io_in_1_acquire_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( io_in_1_acquire_bits_is_builtin_type ),
       .io_in_1_bits_a_type( io_in_1_acquire_bits_a_type ),
       .io_in_1_bits_union( io_in_1_acquire_bits_union ),
       .io_in_1_bits_data( io_in_1_acquire_bits_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_addr_block( io_in_0_acquire_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T56 ),
       .io_in_0_bits_addr_beat( io_in_0_acquire_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( io_in_0_acquire_bits_is_builtin_type ),
       .io_in_0_bits_a_type( io_in_0_acquire_bits_a_type ),
       .io_in_0_bits_union( io_in_0_acquire_bits_union ),
       .io_in_0_bits_data( io_in_0_acquire_bits_data ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( LockingRRArbiter_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( LockingRRArbiter_io_out_bits_a_type ),
       .io_out_bits_union( LockingRRArbiter_io_out_bits_union ),
       .io_out_bits_data( LockingRRArbiter_io_out_bits_data )
       //.io_chosen(  )
  );
endmodule

module L2BroadcastHub(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [127:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data
);

  wire[3:0] T259;
  wire[127:0] T260;
  wire[127:0] T261;
  wire[127:0] T262;
  wire[127:0] T263;
  wire[127:0] T264;
  wire[127:0] T265;
  wire[127:0] T266;
  wire[127:0] T267;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  reg [1:0] rel_data_cnt;
  wire[1:0] T268;
  wire[1:0] T4;
  wire[1:0] T5;
  wire vwbdq_enq;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T269;
  wire[1:0] T270;
  wire[1:0] T271;
  wire T272;
  wire[3:0] T19;
  reg [3:0] sdq_val;
  wire[3:0] T273;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T274;
  wire sdq_enq;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire[3:0] T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T275;
  wire free_sdq;
  wire T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[3:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T276;
  wire T277;
  wire T58;
  wire T59;
  wire[2:0] acquire_idx;
  wire[2:0] T278;
  wire[2:0] T279;
  wire[2:0] T280;
  wire[2:0] T281;
  wire[2:0] T282;
  wire[2:0] T283;
  wire[2:0] T284;
  wire T285;
  wire[7:0] acquireReadys;
  wire[7:0] T61;
  wire[3:0] T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[3:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire[2:0] T296;
  wire[2:0] T297;
  wire[2:0] T298;
  wire T299;
  wire[7:0] acquireMatches;
  wire[7:0] T69;
  wire[3:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire[3:0] T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T76;
  wire T77;
  wire T78;
  wire block_acquires;
  wire T79;
  wire sdq_rdy;
  wire T80;
  wire T81;
  wire[7:0] acquireConflicts;
  wire[7:0] T82;
  wire[3:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[3:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire T93;
  wire T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[3:0] T103;
  wire[3:0] T104;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[3:0] T117;
  wire[3:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire T121;
  wire T122;
  wire[3:0] T123;
  wire[3:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire[3:0] T131;
  wire[3:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[3:0] T146;
  wire[1:0] T147;
  wire[1:0] T148;
  wire T149;
  wire T150;
  wire[3:0] T151;
  wire[3:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[1:0] T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire[3:0] T165;
  wire[3:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[3:0] T173;
  wire[3:0] T174;
  wire[1:0] T175;
  wire[1:0] T176;
  wire T177;
  wire T178;
  wire[3:0] T179;
  wire[3:0] T180;
  wire[1:0] T181;
  wire[1:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[127:0] T187;
  wire[127:0] T188;
  wire[127:0] T189;
  wire[127:0] T190;
  reg [127:0] vwbdq_0;
  wire[127:0] T191;
  wire T192;
  wire T193;
  wire[3:0] T194;
  wire[1:0] T195;
  reg [127:0] vwbdq_1;
  wire[127:0] T196;
  wire T197;
  wire T198;
  wire T199;
  wire[1:0] T200;
  wire[127:0] T201;
  reg [127:0] vwbdq_2;
  wire[127:0] T202;
  wire T203;
  wire T204;
  reg [127:0] vwbdq_3;
  wire[127:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire[127:0] T211;
  wire[127:0] T212;
  reg [127:0] sdq_0;
  wire[127:0] T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[1:0] T217;
  reg [127:0] sdq_1;
  wire[127:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire[1:0] T222;
  wire[127:0] T223;
  reg [127:0] sdq_2;
  wire[127:0] T224;
  wire T225;
  wire T226;
  reg [127:0] sdq_3;
  wire[127:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire[7:0] releaseReadys;
  wire[7:0] T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire[3:0] T238;
  wire[1:0] T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire[2:0] T245;
  wire[2:0] T306;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_probe_valid;
  wire BroadcastVoluntaryReleaseTracker_io_inner_release_ready;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data;
  wire BroadcastVoluntaryReleaseTracker_io_outer_grant_ready;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_match;
  wire BroadcastAcquireTracker_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_finish_ready;
  wire BroadcastAcquireTracker_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_release_ready;
  wire BroadcastAcquireTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_io_outer_grant_ready;
  wire BroadcastAcquireTracker_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_io_has_acquire_match;
  wire BroadcastAcquireTracker_1_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_1_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_finish_ready;
  wire BroadcastAcquireTracker_1_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_release_ready;
  wire BroadcastAcquireTracker_1_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_1_io_outer_grant_ready;
  wire BroadcastAcquireTracker_1_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_1_io_has_acquire_match;
  wire BroadcastAcquireTracker_2_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_2_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_finish_ready;
  wire BroadcastAcquireTracker_2_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_release_ready;
  wire BroadcastAcquireTracker_2_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_2_io_outer_grant_ready;
  wire BroadcastAcquireTracker_2_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_2_io_has_acquire_match;
  wire BroadcastAcquireTracker_3_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_3_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_finish_ready;
  wire BroadcastAcquireTracker_3_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_release_ready;
  wire BroadcastAcquireTracker_3_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_3_io_outer_grant_ready;
  wire BroadcastAcquireTracker_3_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_3_io_has_acquire_match;
  wire BroadcastAcquireTracker_4_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_4_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_4_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_4_io_inner_finish_ready;
  wire BroadcastAcquireTracker_4_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_4_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_4_io_inner_release_ready;
  wire BroadcastAcquireTracker_4_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_4_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_4_io_outer_grant_ready;
  wire BroadcastAcquireTracker_4_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_4_io_has_acquire_match;
  wire BroadcastAcquireTracker_5_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_5_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_5_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_5_io_inner_finish_ready;
  wire BroadcastAcquireTracker_5_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_5_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_5_io_inner_release_ready;
  wire BroadcastAcquireTracker_5_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_5_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_5_io_outer_grant_ready;
  wire BroadcastAcquireTracker_5_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_5_io_has_acquire_match;
  wire BroadcastAcquireTracker_6_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_6_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat;
  wire[5:0] BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_6_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_6_io_inner_finish_ready;
  wire BroadcastAcquireTracker_6_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_6_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_6_io_inner_release_ready;
  wire BroadcastAcquireTracker_6_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block;
  wire[3:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_6_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_6_io_outer_grant_ready;
  wire BroadcastAcquireTracker_6_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_6_io_has_acquire_match;
  wire LockingRRArbiter_io_in_7_ready;
  wire LockingRRArbiter_io_in_6_ready;
  wire LockingRRArbiter_io_in_5_ready;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[5:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[3:0] LockingRRArbiter_io_out_bits_manager_xact_id;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[3:0] LockingRRArbiter_io_out_bits_g_type;
  wire[1:0] LockingRRArbiter_io_out_bits_client_id;
  wire LockingRRArbiter_1_io_in_7_ready;
  wire LockingRRArbiter_1_io_in_6_ready;
  wire LockingRRArbiter_1_io_in_5_ready;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[25:0] LockingRRArbiter_1_io_out_bits_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_p_type;
  wire[1:0] LockingRRArbiter_1_io_out_bits_client_id;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_7_grant_bits_client_xact_id;
  wire outer_arb_io_in_7_grant_bits_manager_xact_id;
  wire outer_arb_io_in_7_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_7_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_7_grant_bits_data;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_6_grant_bits_client_xact_id;
  wire outer_arb_io_in_6_grant_bits_manager_xact_id;
  wire outer_arb_io_in_6_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_6_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_6_grant_bits_data;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_5_grant_bits_client_xact_id;
  wire outer_arb_io_in_5_grant_bits_manager_xact_id;
  wire outer_arb_io_in_5_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_5_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_5_grant_bits_data;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_data;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_data;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_data;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_data;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_data;
  wire outer_arb_io_out_acquire_valid;
  wire[25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire[3:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire[1:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire outer_arb_io_out_acquire_bits_is_builtin_type;
  wire[2:0] outer_arb_io_out_acquire_bits_a_type;
  wire[16:0] outer_arb_io_out_acquire_bits_union;
  wire[3:0] outer_arb_io_out_acquire_bits_data;
  wire outer_arb_io_out_grant_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rel_data_cnt = {1{$random}};
    sdq_val = {1{$random}};
    vwbdq_0 = {4{$random}};
    vwbdq_1 = {4{$random}};
    vwbdq_2 = {4{$random}};
    vwbdq_3 = {4{$random}};
    sdq_0 = {4{$random}};
    sdq_1 = {4{$random}};
    sdq_2 = {4{$random}};
    sdq_3 = {4{$random}};
  end
// synthesis translate_on
`endif

  assign T259 = io_outer_grant_bits_data[2'h3:1'h0];
  assign T260 = {124'h0, BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data};
  assign T261 = {124'h0, BroadcastAcquireTracker_io_inner_grant_bits_data};
  assign T262 = {124'h0, BroadcastAcquireTracker_1_io_inner_grant_bits_data};
  assign T263 = {124'h0, BroadcastAcquireTracker_2_io_inner_grant_bits_data};
  assign T264 = {124'h0, BroadcastAcquireTracker_3_io_inner_grant_bits_data};
  assign T265 = {124'h0, BroadcastAcquireTracker_4_io_inner_grant_bits_data};
  assign T266 = {124'h0, BroadcastAcquireTracker_5_io_inner_grant_bits_data};
  assign T267 = {124'h0, BroadcastAcquireTracker_6_io_inner_grant_bits_data};
  assign T0 = T1;
  assign T1 = {T3, T2};
  assign T2 = 2'h2;
  assign T3 = rel_data_cnt;
  assign T268 = reset ? 2'h0 : T4;
  assign T4 = vwbdq_enq ? T5 : rel_data_cnt;
  assign T5 = rel_data_cnt + 2'h1;
  assign vwbdq_enq = T11 & T6;
  assign T6 = T8 | T7;
  assign T7 = 3'h2 == io_inner_release_bits_r_type;
  assign T8 = T10 | T9;
  assign T9 = 3'h1 == io_inner_release_bits_r_type;
  assign T10 = 3'h0 == io_inner_release_bits_r_type;
  assign T11 = T12 & io_inner_release_bits_voluntary;
  assign T12 = io_inner_release_ready & io_inner_release_valid;
  assign T13 = io_inner_finish_valid & T14;
  assign T14 = io_inner_finish_bits_manager_xact_id == 4'h7;
  assign T15 = T16;
  assign T16 = {T18, T17};
  assign T17 = 2'h0;
  assign T18 = T269;
  assign T269 = T277 ? 1'h0 : T270;
  assign T270 = T276 ? 1'h1 : T271;
  assign T271 = T272 ? 2'h2 : 2'h3;
  assign T272 = T19[2'h2];
  assign T19 = ~ sdq_val;
  assign T273 = reset ? 4'h0 : T20;
  assign T20 = T57 ? T21 : sdq_val;
  assign T21 = T41 | T22;
  assign T22 = T31 & T23;
  assign T23 = 4'h0 - T274;
  assign T274 = {3'h0, sdq_enq};
  assign sdq_enq = T30 & T24;
  assign T24 = io_inner_acquire_bits_is_builtin_type & T25;
  assign T25 = T27 | T26;
  assign T26 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T29 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T30 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T31 = T40 ? 4'h1 : T32;
  assign T32 = T39 ? 4'h2 : T33;
  assign T33 = T38 ? 4'h4 : T34;
  assign T34 = T35 ? 4'h8 : 4'h0;
  assign T35 = T36[2'h3];
  assign T36 = ~ T37;
  assign T37 = sdq_val;
  assign T38 = T36[2'h2];
  assign T39 = T36[1'h1];
  assign T40 = T36[1'h0];
  assign T41 = sdq_val & T42;
  assign T42 = ~ T43;
  assign T43 = T55 & T44;
  assign T44 = 4'h0 - T275;
  assign T275 = {3'h0, free_sdq};
  assign free_sdq = T47 & T45;
  assign T45 = T46 == 2'h0;
  assign T46 = outer_arb_io_out_acquire_bits_data[1'h1:1'h0];
  assign T47 = T54 & T48;
  assign T48 = io_outer_acquire_bits_is_builtin_type & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h4 == io_outer_acquire_bits_a_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T53 = 3'h2 == io_outer_acquire_bits_a_type;
  assign T54 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T55 = 1'h1 << T56;
  assign T56 = outer_arb_io_out_acquire_bits_data[2'h3:2'h2];
  assign T57 = io_outer_acquire_valid | sdq_enq;
  assign T276 = T19[1'h1];
  assign T277 = T19[1'h0];
  assign T58 = T77 & T59;
  assign T59 = acquire_idx == 3'h7;
  assign acquire_idx = T76 ? T292 : T278;
  assign T278 = T291 ? 1'h0 : T279;
  assign T279 = T290 ? 1'h1 : T280;
  assign T280 = T289 ? 2'h2 : T281;
  assign T281 = T288 ? 2'h3 : T282;
  assign T282 = T287 ? 3'h4 : T283;
  assign T283 = T286 ? 3'h5 : T284;
  assign T284 = T285 ? 3'h6 : 3'h7;
  assign T285 = acquireReadys[3'h6];
  assign acquireReadys = T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = {BroadcastAcquireTracker_io_inner_acquire_ready, BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready};
  assign T64 = {BroadcastAcquireTracker_2_io_inner_acquire_ready, BroadcastAcquireTracker_1_io_inner_acquire_ready};
  assign T65 = {T67, T66};
  assign T66 = {BroadcastAcquireTracker_4_io_inner_acquire_ready, BroadcastAcquireTracker_3_io_inner_acquire_ready};
  assign T67 = {BroadcastAcquireTracker_6_io_inner_acquire_ready, BroadcastAcquireTracker_5_io_inner_acquire_ready};
  assign T286 = acquireReadys[3'h5];
  assign T287 = acquireReadys[3'h4];
  assign T288 = acquireReadys[2'h3];
  assign T289 = acquireReadys[2'h2];
  assign T290 = acquireReadys[1'h1];
  assign T291 = acquireReadys[1'h0];
  assign T292 = T305 ? 1'h0 : T293;
  assign T293 = T304 ? 1'h1 : T294;
  assign T294 = T303 ? 2'h2 : T295;
  assign T295 = T302 ? 2'h3 : T296;
  assign T296 = T301 ? 3'h4 : T297;
  assign T297 = T300 ? 3'h5 : T298;
  assign T298 = T299 ? 3'h6 : 3'h7;
  assign T299 = acquireMatches[3'h6];
  assign acquireMatches = T69;
  assign T69 = {T73, T70};
  assign T70 = {T72, T71};
  assign T71 = {BroadcastAcquireTracker_io_has_acquire_match, BroadcastVoluntaryReleaseTracker_io_has_acquire_match};
  assign T72 = {BroadcastAcquireTracker_2_io_has_acquire_match, BroadcastAcquireTracker_1_io_has_acquire_match};
  assign T73 = {T75, T74};
  assign T74 = {BroadcastAcquireTracker_4_io_has_acquire_match, BroadcastAcquireTracker_3_io_has_acquire_match};
  assign T75 = {BroadcastAcquireTracker_6_io_has_acquire_match, BroadcastAcquireTracker_5_io_has_acquire_match};
  assign T300 = acquireMatches[3'h5];
  assign T301 = acquireMatches[3'h4];
  assign T302 = acquireMatches[2'h3];
  assign T303 = acquireMatches[2'h2];
  assign T304 = acquireMatches[1'h1];
  assign T305 = acquireMatches[1'h0];
  assign T76 = acquireMatches != 8'h0;
  assign T77 = io_inner_acquire_valid & T78;
  assign T78 = block_acquires ^ 1'h1;
  assign block_acquires = T81 | T79;
  assign T79 = sdq_rdy ^ 1'h1;
  assign sdq_rdy = T80 ^ 1'h1;
  assign T80 = sdq_val == 4'hf;
  assign T81 = acquireConflicts != 8'h0;
  assign acquireConflicts = T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = {BroadcastAcquireTracker_io_has_acquire_conflict, BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict};
  assign T85 = {BroadcastAcquireTracker_2_io_has_acquire_conflict, BroadcastAcquireTracker_1_io_has_acquire_conflict};
  assign T86 = {T88, T87};
  assign T87 = {BroadcastAcquireTracker_4_io_has_acquire_conflict, BroadcastAcquireTracker_3_io_has_acquire_conflict};
  assign T88 = {BroadcastAcquireTracker_6_io_has_acquire_conflict, BroadcastAcquireTracker_5_io_has_acquire_conflict};
  assign T89 = T90;
  assign T90 = {T92, T91};
  assign T91 = 2'h2;
  assign T92 = rel_data_cnt;
  assign T93 = io_inner_finish_valid & T94;
  assign T94 = io_inner_finish_bits_manager_xact_id == 4'h6;
  assign T95 = T96;
  assign T96 = {T98, T97};
  assign T97 = 2'h0;
  assign T98 = T269;
  assign T99 = T101 & T100;
  assign T100 = acquire_idx == 3'h6;
  assign T101 = io_inner_acquire_valid & T102;
  assign T102 = block_acquires ^ 1'h1;
  assign T103 = T104;
  assign T104 = {T106, T105};
  assign T105 = 2'h2;
  assign T106 = rel_data_cnt;
  assign T107 = io_inner_finish_valid & T108;
  assign T108 = io_inner_finish_bits_manager_xact_id == 4'h5;
  assign T109 = T110;
  assign T110 = {T112, T111};
  assign T111 = 2'h0;
  assign T112 = T269;
  assign T113 = T115 & T114;
  assign T114 = acquire_idx == 3'h5;
  assign T115 = io_inner_acquire_valid & T116;
  assign T116 = block_acquires ^ 1'h1;
  assign T117 = T118;
  assign T118 = {T120, T119};
  assign T119 = 2'h2;
  assign T120 = rel_data_cnt;
  assign T121 = io_inner_finish_valid & T122;
  assign T122 = io_inner_finish_bits_manager_xact_id == 4'h4;
  assign T123 = T124;
  assign T124 = {T126, T125};
  assign T125 = 2'h0;
  assign T126 = T269;
  assign T127 = T129 & T128;
  assign T128 = acquire_idx == 3'h4;
  assign T129 = io_inner_acquire_valid & T130;
  assign T130 = block_acquires ^ 1'h1;
  assign T131 = T132;
  assign T132 = {T134, T133};
  assign T133 = 2'h2;
  assign T134 = rel_data_cnt;
  assign T135 = io_inner_finish_valid & T136;
  assign T136 = io_inner_finish_bits_manager_xact_id == 4'h3;
  assign T137 = T138;
  assign T138 = {T140, T139};
  assign T139 = 2'h0;
  assign T140 = T269;
  assign T141 = T143 & T142;
  assign T142 = acquire_idx == 3'h3;
  assign T143 = io_inner_acquire_valid & T144;
  assign T144 = block_acquires ^ 1'h1;
  assign T145 = T146;
  assign T146 = {T148, T147};
  assign T147 = 2'h2;
  assign T148 = rel_data_cnt;
  assign T149 = io_inner_finish_valid & T150;
  assign T150 = io_inner_finish_bits_manager_xact_id == 4'h2;
  assign T151 = T152;
  assign T152 = {T154, T153};
  assign T153 = 2'h0;
  assign T154 = T269;
  assign T155 = T157 & T156;
  assign T156 = acquire_idx == 3'h2;
  assign T157 = io_inner_acquire_valid & T158;
  assign T158 = block_acquires ^ 1'h1;
  assign T159 = T160;
  assign T160 = {T162, T161};
  assign T161 = 2'h2;
  assign T162 = rel_data_cnt;
  assign T163 = io_inner_finish_valid & T164;
  assign T164 = io_inner_finish_bits_manager_xact_id == 4'h1;
  assign T165 = T166;
  assign T166 = {T168, T167};
  assign T167 = 2'h0;
  assign T168 = T269;
  assign T169 = T171 & T170;
  assign T170 = acquire_idx == 3'h1;
  assign T171 = io_inner_acquire_valid & T172;
  assign T172 = block_acquires ^ 1'h1;
  assign T173 = T174;
  assign T174 = {T176, T175};
  assign T175 = 2'h1;
  assign T176 = rel_data_cnt;
  assign T177 = io_inner_finish_valid & T178;
  assign T178 = io_inner_finish_bits_manager_xact_id == 4'h0;
  assign T179 = T180;
  assign T180 = {T182, T181};
  assign T181 = 2'h0;
  assign T182 = T269;
  assign T183 = T185 & T184;
  assign T184 = acquire_idx == 3'h0;
  assign T185 = io_inner_acquire_valid & T186;
  assign T186 = block_acquires ^ 1'h1;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_data = T187;
  assign T187 = T232 ? T211 : T188;
  assign T188 = T210 ? T189 : io_inner_release_bits_data;
  assign T189 = T209 ? T201 : T190;
  assign T190 = T199 ? vwbdq_1 : vwbdq_0;
  assign T191 = T192 ? io_inner_release_bits_data : vwbdq_0;
  assign T192 = vwbdq_enq & T193;
  assign T193 = T194[1'h0];
  assign T194 = 1'h1 << T195;
  assign T195 = rel_data_cnt;
  assign T196 = T197 ? io_inner_release_bits_data : vwbdq_1;
  assign T197 = vwbdq_enq & T198;
  assign T198 = T194[1'h1];
  assign T199 = T200[1'h0];
  assign T200 = T56;
  assign T201 = T208 ? vwbdq_3 : vwbdq_2;
  assign T202 = T203 ? io_inner_release_bits_data : vwbdq_2;
  assign T203 = vwbdq_enq & T204;
  assign T204 = T194[2'h2];
  assign T205 = T206 ? io_inner_release_bits_data : vwbdq_3;
  assign T206 = vwbdq_enq & T207;
  assign T207 = T194[2'h3];
  assign T208 = T200[1'h0];
  assign T209 = T200[1'h1];
  assign T210 = T46 == 2'h1;
  assign T211 = T231 ? T223 : T212;
  assign T212 = T221 ? sdq_1 : sdq_0;
  assign T213 = T214 ? io_inner_acquire_bits_data : sdq_0;
  assign T214 = sdq_enq & T215;
  assign T215 = T216[1'h0];
  assign T216 = 1'h1 << T217;
  assign T217 = T269;
  assign T218 = T219 ? io_inner_acquire_bits_data : sdq_1;
  assign T219 = sdq_enq & T220;
  assign T220 = T216[1'h1];
  assign T221 = T222[1'h0];
  assign T222 = T56;
  assign T223 = T230 ? sdq_3 : sdq_2;
  assign T224 = T225 ? io_inner_acquire_bits_data : sdq_2;
  assign T225 = sdq_enq & T226;
  assign T226 = T216[2'h2];
  assign T227 = T228 ? io_inner_acquire_bits_data : sdq_3;
  assign T228 = sdq_enq & T229;
  assign T229 = T216[2'h3];
  assign T230 = T222[1'h0];
  assign T231 = T222[1'h1];
  assign T232 = T46 == 2'h0;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T233;
  assign T233 = releaseReadys != 8'h0;
  assign releaseReadys = T234;
  assign T234 = {T238, T235};
  assign T235 = {T237, T236};
  assign T236 = {BroadcastAcquireTracker_io_inner_release_ready, BroadcastVoluntaryReleaseTracker_io_inner_release_ready};
  assign T237 = {BroadcastAcquireTracker_2_io_inner_release_ready, BroadcastAcquireTracker_1_io_inner_release_ready};
  assign T238 = {T240, T239};
  assign T239 = {BroadcastAcquireTracker_4_io_inner_release_ready, BroadcastAcquireTracker_3_io_inner_release_ready};
  assign T240 = {BroadcastAcquireTracker_6_io_inner_release_ready, BroadcastAcquireTracker_5_io_inner_release_ready};
  assign io_inner_probe_bits_client_id = LockingRRArbiter_1_io_out_bits_client_id;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_1_io_out_bits_p_type;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_1_io_out_bits_addr_block;
  assign io_inner_probe_valid = LockingRRArbiter_1_io_out_valid;
  assign io_inner_finish_ready = T241;
  assign T241 = T255 ? T249 : T242;
  assign T242 = T248 ? T246 : T243;
  assign T243 = T244 ? BroadcastAcquireTracker_io_inner_finish_ready : BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  assign T244 = T245[1'h0];
  assign T245 = T306;
  assign T306 = io_inner_finish_bits_manager_xact_id[2'h2:1'h0];
  assign T246 = T247 ? BroadcastAcquireTracker_2_io_inner_finish_ready : BroadcastAcquireTracker_1_io_inner_finish_ready;
  assign T247 = T245[1'h0];
  assign T248 = T245[1'h1];
  assign T249 = T254 ? T252 : T250;
  assign T250 = T251 ? BroadcastAcquireTracker_4_io_inner_finish_ready : BroadcastAcquireTracker_3_io_inner_finish_ready;
  assign T251 = T245[1'h0];
  assign T252 = T253 ? BroadcastAcquireTracker_6_io_inner_finish_ready : BroadcastAcquireTracker_5_io_inner_finish_ready;
  assign T253 = T245[1'h0];
  assign T254 = T245[1'h1];
  assign T255 = T245[2'h2];
  assign io_inner_grant_bits_client_id = LockingRRArbiter_io_out_bits_client_id;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_io_out_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = LockingRRArbiter_io_out_valid;
  assign io_inner_acquire_ready = T256;
  assign T256 = T258 & T257;
  assign T257 = block_acquires ^ 1'h1;
  assign T258 = acquireReadys != 8'h0;
  BroadcastVoluntaryReleaseTracker BroadcastVoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T183 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T179 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_0_ready ),
       .io_inner_grant_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastVoluntaryReleaseTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T177 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_inner_probe_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_addr_block(  )
       //.io_inner_probe_bits_p_type(  )
       //.io_inner_probe_bits_client_id(  )
       .io_inner_release_ready( BroadcastVoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T173 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastVoluntaryReleaseTracker_io_has_acquire_match )
  );
  BroadcastAcquireTracker_0 BroadcastAcquireTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T169 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T165 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_1_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T163 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T159 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_io_has_acquire_match )
  );
  BroadcastAcquireTracker_1 BroadcastAcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T155 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T151 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_2_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_1_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_1_io_inner_finish_ready ),
       .io_inner_finish_valid( T149 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T145 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_1_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_1_io_has_acquire_match )
  );
  BroadcastAcquireTracker_2 BroadcastAcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T141 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T137 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_3_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_2_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_2_io_inner_finish_ready ),
       .io_inner_finish_valid( T135 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T131 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_2_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_2_io_has_acquire_match )
  );
  BroadcastAcquireTracker_3 BroadcastAcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T127 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T123 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_4_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_3_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_3_io_inner_finish_ready ),
       .io_inner_finish_valid( T121 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T117 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_3_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_3_io_has_acquire_match )
  );
  BroadcastAcquireTracker_4 BroadcastAcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T113 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T109 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_5_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_4_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_4_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_4_io_inner_finish_ready ),
       .io_inner_finish_valid( T107 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_5_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_4_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_4_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T103 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_4_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_4_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_5_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_5_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_5_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_5_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_5_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_5_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_4_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_4_io_has_acquire_match )
  );
  BroadcastAcquireTracker_5 BroadcastAcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T99 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T95 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_6_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_5_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_5_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_5_io_inner_finish_ready ),
       .io_inner_finish_valid( T93 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_6_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_5_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_5_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T89 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_5_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_5_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_6_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_6_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_6_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_6_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_6_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_6_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_5_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_5_io_has_acquire_match )
  );
  BroadcastAcquireTracker_6 BroadcastAcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T58 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T15 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_7_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_6_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_6_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_6_io_inner_finish_ready ),
       .io_inner_finish_valid( T13 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_7_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_6_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_6_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( io_inner_release_valid ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T0 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_6_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_6_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_7_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_7_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_7_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_7_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_7_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_7_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_6_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_6_io_has_acquire_match )
  );
  LockingRRArbiter_2 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_io_in_7_ready ),
       .io_in_7_valid( BroadcastAcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_addr_beat( BroadcastAcquireTracker_6_io_inner_grant_bits_addr_beat ),
       .io_in_7_bits_client_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_xact_id ),
       .io_in_7_bits_manager_xact_id( BroadcastAcquireTracker_6_io_inner_grant_bits_manager_xact_id ),
       .io_in_7_bits_is_builtin_type( BroadcastAcquireTracker_6_io_inner_grant_bits_is_builtin_type ),
       .io_in_7_bits_g_type( BroadcastAcquireTracker_6_io_inner_grant_bits_g_type ),
       .io_in_7_bits_data( T267 ),
       .io_in_7_bits_client_id( BroadcastAcquireTracker_6_io_inner_grant_bits_client_id ),
       .io_in_6_ready( LockingRRArbiter_io_in_6_ready ),
       .io_in_6_valid( BroadcastAcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_addr_beat( BroadcastAcquireTracker_5_io_inner_grant_bits_addr_beat ),
       .io_in_6_bits_client_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_xact_id ),
       .io_in_6_bits_manager_xact_id( BroadcastAcquireTracker_5_io_inner_grant_bits_manager_xact_id ),
       .io_in_6_bits_is_builtin_type( BroadcastAcquireTracker_5_io_inner_grant_bits_is_builtin_type ),
       .io_in_6_bits_g_type( BroadcastAcquireTracker_5_io_inner_grant_bits_g_type ),
       .io_in_6_bits_data( T266 ),
       .io_in_6_bits_client_id( BroadcastAcquireTracker_5_io_inner_grant_bits_client_id ),
       .io_in_5_ready( LockingRRArbiter_io_in_5_ready ),
       .io_in_5_valid( BroadcastAcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_addr_beat( BroadcastAcquireTracker_4_io_inner_grant_bits_addr_beat ),
       .io_in_5_bits_client_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_xact_id ),
       .io_in_5_bits_manager_xact_id( BroadcastAcquireTracker_4_io_inner_grant_bits_manager_xact_id ),
       .io_in_5_bits_is_builtin_type( BroadcastAcquireTracker_4_io_inner_grant_bits_is_builtin_type ),
       .io_in_5_bits_g_type( BroadcastAcquireTracker_4_io_inner_grant_bits_g_type ),
       .io_in_5_bits_data( T265 ),
       .io_in_5_bits_client_id( BroadcastAcquireTracker_4_io_inner_grant_bits_client_id ),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_in_4_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_in_4_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_in_4_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_in_4_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_in_4_bits_data( T264 ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_in_3_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_in_3_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_in_3_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_in_3_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_in_3_bits_data( T263 ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_in_2_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_in_2_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_in_2_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_in_2_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_in_2_bits_data( T262 ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_in_1_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_in_1_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_1_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_1_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_1_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_in_1_bits_data( T261 ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_in_0_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_0_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_0_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_0_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_in_0_bits_data( T260 ),
       .io_in_0_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( LockingRRArbiter_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( LockingRRArbiter_io_out_bits_g_type ),
       //.io_out_bits_data(  )
       .io_out_bits_client_id( LockingRRArbiter_io_out_bits_client_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_1_io_in_7_ready ),
       .io_in_7_valid( BroadcastAcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_addr_block( BroadcastAcquireTracker_6_io_inner_probe_bits_addr_block ),
       .io_in_7_bits_p_type( BroadcastAcquireTracker_6_io_inner_probe_bits_p_type ),
       .io_in_7_bits_client_id( BroadcastAcquireTracker_6_io_inner_probe_bits_client_id ),
       .io_in_6_ready( LockingRRArbiter_1_io_in_6_ready ),
       .io_in_6_valid( BroadcastAcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_addr_block( BroadcastAcquireTracker_5_io_inner_probe_bits_addr_block ),
       .io_in_6_bits_p_type( BroadcastAcquireTracker_5_io_inner_probe_bits_p_type ),
       .io_in_6_bits_client_id( BroadcastAcquireTracker_5_io_inner_probe_bits_client_id ),
       .io_in_5_ready( LockingRRArbiter_1_io_in_5_ready ),
       .io_in_5_valid( BroadcastAcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_addr_block( BroadcastAcquireTracker_4_io_inner_probe_bits_addr_block ),
       .io_in_5_bits_p_type( BroadcastAcquireTracker_4_io_inner_probe_bits_p_type ),
       .io_in_5_bits_client_id( BroadcastAcquireTracker_4_io_inner_probe_bits_client_id ),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_in_4_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_in_3_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_in_2_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_in_1_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_in_1_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_addr_block(  )
       //.io_in_0_bits_p_type(  )
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_1_io_out_bits_addr_block ),
       .io_out_bits_p_type( LockingRRArbiter_1_io_out_bits_p_type ),
       .io_out_bits_client_id( LockingRRArbiter_1_io_out_bits_client_id )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign LockingRRArbiter_1.io_in_0_bits_addr_block = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_p_type = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  ClientUncachedTileLinkIOArbiter outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( BroadcastAcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_addr_block( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_block ),
       .io_in_7_acquire_bits_client_xact_id( BroadcastAcquireTracker_6_io_outer_acquire_bits_client_xact_id ),
       .io_in_7_acquire_bits_addr_beat( BroadcastAcquireTracker_6_io_outer_acquire_bits_addr_beat ),
       .io_in_7_acquire_bits_is_builtin_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_is_builtin_type ),
       .io_in_7_acquire_bits_a_type( BroadcastAcquireTracker_6_io_outer_acquire_bits_a_type ),
       .io_in_7_acquire_bits_union( BroadcastAcquireTracker_6_io_outer_acquire_bits_union ),
       .io_in_7_acquire_bits_data( BroadcastAcquireTracker_6_io_outer_acquire_bits_data ),
       .io_in_7_grant_ready( BroadcastAcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_addr_beat( outer_arb_io_in_7_grant_bits_addr_beat ),
       .io_in_7_grant_bits_client_xact_id( outer_arb_io_in_7_grant_bits_client_xact_id ),
       .io_in_7_grant_bits_manager_xact_id( outer_arb_io_in_7_grant_bits_manager_xact_id ),
       .io_in_7_grant_bits_is_builtin_type( outer_arb_io_in_7_grant_bits_is_builtin_type ),
       .io_in_7_grant_bits_g_type( outer_arb_io_in_7_grant_bits_g_type ),
       .io_in_7_grant_bits_data( outer_arb_io_in_7_grant_bits_data ),
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( BroadcastAcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_addr_block( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_block ),
       .io_in_6_acquire_bits_client_xact_id( BroadcastAcquireTracker_5_io_outer_acquire_bits_client_xact_id ),
       .io_in_6_acquire_bits_addr_beat( BroadcastAcquireTracker_5_io_outer_acquire_bits_addr_beat ),
       .io_in_6_acquire_bits_is_builtin_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_is_builtin_type ),
       .io_in_6_acquire_bits_a_type( BroadcastAcquireTracker_5_io_outer_acquire_bits_a_type ),
       .io_in_6_acquire_bits_union( BroadcastAcquireTracker_5_io_outer_acquire_bits_union ),
       .io_in_6_acquire_bits_data( BroadcastAcquireTracker_5_io_outer_acquire_bits_data ),
       .io_in_6_grant_ready( BroadcastAcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_addr_beat( outer_arb_io_in_6_grant_bits_addr_beat ),
       .io_in_6_grant_bits_client_xact_id( outer_arb_io_in_6_grant_bits_client_xact_id ),
       .io_in_6_grant_bits_manager_xact_id( outer_arb_io_in_6_grant_bits_manager_xact_id ),
       .io_in_6_grant_bits_is_builtin_type( outer_arb_io_in_6_grant_bits_is_builtin_type ),
       .io_in_6_grant_bits_g_type( outer_arb_io_in_6_grant_bits_g_type ),
       .io_in_6_grant_bits_data( outer_arb_io_in_6_grant_bits_data ),
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( BroadcastAcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_addr_block( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_block ),
       .io_in_5_acquire_bits_client_xact_id( BroadcastAcquireTracker_4_io_outer_acquire_bits_client_xact_id ),
       .io_in_5_acquire_bits_addr_beat( BroadcastAcquireTracker_4_io_outer_acquire_bits_addr_beat ),
       .io_in_5_acquire_bits_is_builtin_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_is_builtin_type ),
       .io_in_5_acquire_bits_a_type( BroadcastAcquireTracker_4_io_outer_acquire_bits_a_type ),
       .io_in_5_acquire_bits_union( BroadcastAcquireTracker_4_io_outer_acquire_bits_union ),
       .io_in_5_acquire_bits_data( BroadcastAcquireTracker_4_io_outer_acquire_bits_data ),
       .io_in_5_grant_ready( BroadcastAcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_addr_beat( outer_arb_io_in_5_grant_bits_addr_beat ),
       .io_in_5_grant_bits_client_xact_id( outer_arb_io_in_5_grant_bits_client_xact_id ),
       .io_in_5_grant_bits_manager_xact_id( outer_arb_io_in_5_grant_bits_manager_xact_id ),
       .io_in_5_grant_bits_is_builtin_type( outer_arb_io_in_5_grant_bits_is_builtin_type ),
       .io_in_5_grant_bits_g_type( outer_arb_io_in_5_grant_bits_g_type ),
       .io_in_5_grant_bits_data( outer_arb_io_in_5_grant_bits_data ),
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_in_4_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_in_4_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_in_4_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_in_4_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_in_4_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_in_4_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_in_4_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_in_4_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_in_4_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_in_4_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_in_4_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_in_4_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_in_3_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_in_3_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_in_3_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_in_3_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_in_3_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_in_3_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_in_3_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_in_3_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_in_3_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_in_3_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_in_3_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_in_3_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_in_2_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_in_2_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_in_2_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_in_2_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_in_2_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_in_2_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_in_2_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_in_2_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_in_2_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_in_2_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_in_2_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_in_2_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_in_1_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_1_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_1_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_1_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_in_1_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_in_1_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_in_1_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_in_1_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_in_1_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_in_1_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_in_1_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_in_1_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_in_0_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_0_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_0_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_0_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_in_0_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_in_0_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_in_0_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_in_0_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_in_0_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_in_0_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_in_0_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_in_0_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( outer_arb_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( outer_arb_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( outer_arb_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( outer_arb_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( outer_arb_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( outer_arb_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( outer_arb_io_out_acquire_bits_data ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_addr_beat( io_outer_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( io_outer_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( io_outer_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( io_outer_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( io_outer_grant_bits_g_type ),
       .io_out_grant_bits_data( T259 )
  );

  always @(posedge clk) begin
    if(reset) begin
      rel_data_cnt <= 2'h0;
    end else if(vwbdq_enq) begin
      rel_data_cnt <= T5;
    end
    if(reset) begin
      sdq_val <= 4'h0;
    end else if(T57) begin
      sdq_val <= T21;
    end
    if(T192) begin
      vwbdq_0 <= io_inner_release_bits_data;
    end
    if(T197) begin
      vwbdq_1 <= io_inner_release_bits_data;
    end
    if(T203) begin
      vwbdq_2 <= io_inner_release_bits_data;
    end
    if(T206) begin
      vwbdq_3 <= io_inner_release_bits_data;
    end
    if(T214) begin
      sdq_0 <= io_inner_acquire_bits_data;
    end
    if(T219) begin
      sdq_1 <= io_inner_acquire_bits_data;
    end
    if(T225) begin
      sdq_2 <= io_inner_acquire_bits_data;
    end
    if(T228) begin
      sdq_3 <= io_inner_acquire_bits_data;
    end
  end
endmodule

module MMIOTileLinkManager(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [5:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[5:0] io_inner_grant_bits_client_xact_id,
    output[3:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [3:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[25:0] io_inner_probe_bits_addr_block
    //output[1:0] io_inner_probe_bits_p_type
    //output[1:0] io_inner_probe_bits_client_id
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [5:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [127:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    //input  io_incoherent_0
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data
);

  wire[3:0] outer_xact_id;
  wire[3:0] T134;
  wire[3:0] T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire[8:0] T0;
  reg [8:0] xact_pending;
  wire[8:0] T143;
  wire[15:0] T144;
  wire[15:0] T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[15:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[15:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire[15:0] T23;
  wire T24;
  wire[15:0] T25;
  wire[15:0] T26;
  wire[15:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[15:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg [3:0] xact_id_reg;
  wire[3:0] T35;
  wire multibeat_start;
  wire T36;
  wire multibeat_fire;
  wire T37;
  wire T38;
  wire T39;
  reg  xact_multibeat;
  wire T153;
  wire T40;
  wire T41;
  wire multibeat_end;
  wire T42;
  wire T43;
  wire xact_free;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  reg [1:0] xact_buffer_0_client_id;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire[15:0] T53;
  wire[3:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  reg [1:0] xact_buffer_1_client_id;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[1:0] T67;
  reg [1:0] xact_buffer_2_client_id;
  wire[1:0] T68;
  wire T69;
  wire T70;
  reg [1:0] xact_buffer_3_client_id;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[1:0] T76;
  wire[1:0] T77;
  reg [1:0] xact_buffer_4_client_id;
  wire[1:0] T78;
  wire T79;
  wire T80;
  reg [1:0] xact_buffer_5_client_id;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire[1:0] T85;
  reg [1:0] xact_buffer_6_client_id;
  wire[1:0] T86;
  wire T87;
  wire T88;
  reg [1:0] xact_buffer_7_client_id;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  reg [1:0] xact_buffer_8_client_id;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[5:0] T99;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  reg [5:0] xact_buffer_0_client_xact_id;
  wire[5:0] T103;
  wire T104;
  reg [5:0] xact_buffer_1_client_xact_id;
  wire[5:0] T105;
  wire T106;
  wire T107;
  wire[5:0] T108;
  reg [5:0] xact_buffer_2_client_xact_id;
  wire[5:0] T109;
  wire T110;
  reg [5:0] xact_buffer_3_client_xact_id;
  wire[5:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[5:0] T115;
  wire[5:0] T116;
  reg [5:0] xact_buffer_4_client_xact_id;
  wire[5:0] T117;
  wire T118;
  reg [5:0] xact_buffer_5_client_xact_id;
  wire[5:0] T119;
  wire T120;
  wire T121;
  wire[5:0] T122;
  reg [5:0] xact_buffer_6_client_xact_id;
  wire[5:0] T123;
  wire T124;
  reg [5:0] xact_buffer_7_client_xact_id;
  wire[5:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  reg [5:0] xact_buffer_8_client_xact_id;
  wire[5:0] T130;
  wire T131;
  wire T132;
  wire T133;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    xact_pending = {1{$random}};
    xact_id_reg = {1{$random}};
    xact_multibeat = {1{$random}};
    xact_buffer_0_client_id = {1{$random}};
    xact_buffer_1_client_id = {1{$random}};
    xact_buffer_2_client_id = {1{$random}};
    xact_buffer_3_client_id = {1{$random}};
    xact_buffer_4_client_id = {1{$random}};
    xact_buffer_5_client_id = {1{$random}};
    xact_buffer_6_client_id = {1{$random}};
    xact_buffer_7_client_id = {1{$random}};
    xact_buffer_8_client_id = {1{$random}};
    xact_buffer_0_client_xact_id = {1{$random}};
    xact_buffer_1_client_xact_id = {1{$random}};
    xact_buffer_2_client_xact_id = {1{$random}};
    xact_buffer_3_client_xact_id = {1{$random}};
    xact_buffer_4_client_xact_id = {1{$random}};
    xact_buffer_5_client_xact_id = {1{$random}};
    xact_buffer_6_client_xact_id = {1{$random}};
    xact_buffer_7_client_xact_id = {1{$random}};
    xact_buffer_8_client_xact_id = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_inner_probe_bits_client_id = {1{$random}};
//  assign io_inner_probe_bits_p_type = {1{$random}};
//  assign io_inner_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : T134;
  assign T134 = T152 ? 1'h0 : T135;
  assign T135 = T151 ? 1'h1 : T136;
  assign T136 = T150 ? 2'h2 : T137;
  assign T137 = T149 ? 2'h3 : T138;
  assign T138 = T148 ? 3'h4 : T139;
  assign T139 = T147 ? 3'h5 : T140;
  assign T140 = T146 ? 3'h6 : T141;
  assign T141 = T142 ? 3'h7 : 4'h8;
  assign T142 = T0[3'h7];
  assign T0 = ~ xact_pending;
  assign T143 = T144[4'h8:1'h0];
  assign T144 = reset ? 16'h0 : T1;
  assign T1 = T20 & T2;
  assign T2 = ~ T3;
  assign T3 = T5 ? T4 : 16'h0;
  assign T4 = 1'h1 << io_inner_grant_bits_manager_xact_id;
  assign T5 = T10 & T6;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_inner_grant_bits_is_builtin_type & T9;
  assign T9 = io_inner_grant_bits_g_type == 4'h0;
  assign T10 = T19 & T11;
  assign T11 = T13 | T12;
  assign T12 = io_inner_grant_bits_addr_beat == 2'h3;
  assign T13 = T14 ^ 1'h1;
  assign T14 = io_inner_grant_bits_is_builtin_type ? T18 : T15;
  assign T15 = T17 | T16;
  assign T16 = 4'h1 == io_inner_grant_bits_g_type;
  assign T17 = 4'h0 == io_inner_grant_bits_g_type;
  assign T18 = 4'h5 == io_inner_grant_bits_g_type;
  assign T19 = io_inner_grant_ready & io_inner_grant_valid;
  assign T20 = T25 & T21;
  assign T21 = ~ T22;
  assign T22 = T24 ? T23 : 16'h0;
  assign T23 = 1'h1 << io_inner_finish_bits_manager_xact_id;
  assign T24 = io_inner_finish_ready & io_inner_finish_valid;
  assign T25 = T145 | T26;
  assign T26 = T28 ? T27 : 16'h0;
  assign T27 = 1'h1 << io_outer_acquire_bits_client_xact_id;
  assign T28 = T34 & T29;
  assign T29 = T31 | T30;
  assign T30 = io_outer_acquire_bits_addr_beat == 2'h3;
  assign T31 = T32 ^ 1'h1;
  assign T32 = io_outer_acquire_bits_is_builtin_type & T33;
  assign T33 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T34 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T145 = {7'h0, xact_pending};
  assign T146 = T0[3'h6];
  assign T147 = T0[3'h5];
  assign T148 = T0[3'h4];
  assign T149 = T0[2'h3];
  assign T150 = T0[2'h2];
  assign T151 = T0[1'h1];
  assign T152 = T0[1'h0];
  assign T35 = multibeat_start ? T134 : xact_id_reg;
  assign multibeat_start = multibeat_fire & T36;
  assign T36 = io_outer_acquire_bits_addr_beat == 2'h0;
  assign multibeat_fire = T39 & T37;
  assign T37 = io_outer_acquire_bits_is_builtin_type & T38;
  assign T38 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T39 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T153 = reset ? 1'h0 : T40;
  assign T40 = multibeat_end ? 1'h0 : T41;
  assign T41 = multibeat_start ? 1'h1 : xact_multibeat;
  assign multibeat_end = multibeat_fire & T42;
  assign T42 = io_outer_acquire_bits_addr_beat == 2'h3;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_valid = T43;
  assign T43 = io_inner_acquire_valid & xact_free;
  assign xact_free = T44 ^ 1'h1;
  assign T44 = xact_pending == 9'h1ff;
  assign io_inner_release_ready = 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = T45;
  assign T45 = xact_pending[io_inner_finish_bits_manager_xact_id];
  assign io_inner_grant_bits_client_id = T46;
  assign T46 = T98 ? xact_buffer_8_client_id : T47;
  assign T47 = T94 ? T76 : T48;
  assign T48 = T75 ? T67 : T49;
  assign T49 = T65 ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign T50 = T51 ? io_inner_acquire_bits_client_id : xact_buffer_0_client_id;
  assign T51 = T55 & T52;
  assign T52 = T53[1'h0];
  assign T53 = 1'h1 << T54;
  assign T54 = outer_xact_id;
  assign T55 = T61 & T56;
  assign T56 = T58 | T57;
  assign T57 = io_outer_acquire_bits_addr_beat == 2'h3;
  assign T58 = T59 ^ 1'h1;
  assign T59 = io_outer_acquire_bits_is_builtin_type & T60;
  assign T60 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T61 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T62 = T63 ? io_inner_acquire_bits_client_id : xact_buffer_1_client_id;
  assign T63 = T55 & T64;
  assign T64 = T53[1'h1];
  assign T65 = T66[1'h0];
  assign T66 = io_outer_grant_bits_client_xact_id;
  assign T67 = T74 ? xact_buffer_3_client_id : xact_buffer_2_client_id;
  assign T68 = T69 ? io_inner_acquire_bits_client_id : xact_buffer_2_client_id;
  assign T69 = T55 & T70;
  assign T70 = T53[2'h2];
  assign T71 = T72 ? io_inner_acquire_bits_client_id : xact_buffer_3_client_id;
  assign T72 = T55 & T73;
  assign T73 = T53[2'h3];
  assign T74 = T66[1'h0];
  assign T75 = T66[1'h1];
  assign T76 = T93 ? T85 : T77;
  assign T77 = T84 ? xact_buffer_5_client_id : xact_buffer_4_client_id;
  assign T78 = T79 ? io_inner_acquire_bits_client_id : xact_buffer_4_client_id;
  assign T79 = T55 & T80;
  assign T80 = T53[3'h4];
  assign T81 = T82 ? io_inner_acquire_bits_client_id : xact_buffer_5_client_id;
  assign T82 = T55 & T83;
  assign T83 = T53[3'h5];
  assign T84 = T66[1'h0];
  assign T85 = T92 ? xact_buffer_7_client_id : xact_buffer_6_client_id;
  assign T86 = T87 ? io_inner_acquire_bits_client_id : xact_buffer_6_client_id;
  assign T87 = T55 & T88;
  assign T88 = T53[3'h6];
  assign T89 = T90 ? io_inner_acquire_bits_client_id : xact_buffer_7_client_id;
  assign T90 = T55 & T91;
  assign T91 = T53[3'h7];
  assign T92 = T66[1'h0];
  assign T93 = T66[1'h1];
  assign T94 = T66[2'h2];
  assign T95 = T96 ? io_inner_acquire_bits_client_id : xact_buffer_8_client_id;
  assign T96 = T55 & T97;
  assign T97 = T53[4'h8];
  assign T98 = T66[2'h3];
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_client_xact_id = T99;
  assign T99 = T132 ? xact_buffer_8_client_xact_id : T100;
  assign T100 = T129 ? T115 : T101;
  assign T101 = T114 ? T108 : T102;
  assign T102 = T107 ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign T103 = T104 ? io_inner_acquire_bits_client_xact_id : xact_buffer_0_client_xact_id;
  assign T104 = T55 & T52;
  assign T105 = T106 ? io_inner_acquire_bits_client_xact_id : xact_buffer_1_client_xact_id;
  assign T106 = T55 & T64;
  assign T107 = T66[1'h0];
  assign T108 = T113 ? xact_buffer_3_client_xact_id : xact_buffer_2_client_xact_id;
  assign T109 = T110 ? io_inner_acquire_bits_client_xact_id : xact_buffer_2_client_xact_id;
  assign T110 = T55 & T70;
  assign T111 = T112 ? io_inner_acquire_bits_client_xact_id : xact_buffer_3_client_xact_id;
  assign T112 = T55 & T73;
  assign T113 = T66[1'h0];
  assign T114 = T66[1'h1];
  assign T115 = T128 ? T122 : T116;
  assign T116 = T121 ? xact_buffer_5_client_xact_id : xact_buffer_4_client_xact_id;
  assign T117 = T118 ? io_inner_acquire_bits_client_xact_id : xact_buffer_4_client_xact_id;
  assign T118 = T55 & T80;
  assign T119 = T120 ? io_inner_acquire_bits_client_xact_id : xact_buffer_5_client_xact_id;
  assign T120 = T55 & T83;
  assign T121 = T66[1'h0];
  assign T122 = T127 ? xact_buffer_7_client_xact_id : xact_buffer_6_client_xact_id;
  assign T123 = T124 ? io_inner_acquire_bits_client_xact_id : xact_buffer_6_client_xact_id;
  assign T124 = T55 & T88;
  assign T125 = T126 ? io_inner_acquire_bits_client_xact_id : xact_buffer_7_client_xact_id;
  assign T126 = T55 & T91;
  assign T127 = T66[1'h0];
  assign T128 = T66[1'h1];
  assign T129 = T66[2'h2];
  assign T130 = T131 ? io_inner_acquire_bits_client_xact_id : xact_buffer_8_client_xact_id;
  assign T131 = T55 & T97;
  assign T132 = T66[2'h3];
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_acquire_ready = T133;
  assign T133 = io_outer_acquire_ready & xact_free;

  always @(posedge clk) begin
    xact_pending <= T143;
    if(multibeat_start) begin
      xact_id_reg <= T134;
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else if(multibeat_end) begin
      xact_multibeat <= 1'h0;
    end else if(multibeat_start) begin
      xact_multibeat <= 1'h1;
    end
    if(T51) begin
      xact_buffer_0_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T63) begin
      xact_buffer_1_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T69) begin
      xact_buffer_2_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T72) begin
      xact_buffer_3_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T79) begin
      xact_buffer_4_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T82) begin
      xact_buffer_5_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T87) begin
      xact_buffer_6_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T90) begin
      xact_buffer_7_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T96) begin
      xact_buffer_8_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T104) begin
      xact_buffer_0_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T106) begin
      xact_buffer_1_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T110) begin
      xact_buffer_2_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T112) begin
      xact_buffer_3_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T118) begin
      xact_buffer_4_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T120) begin
      xact_buffer_5_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T124) begin
      xact_buffer_6_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T126) begin
      xact_buffer_7_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(T131) begin
      xact_buffer_8_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_len,
    input [2:0] io_enq_bits_size,
    input [1:0] io_enq_bits_burst,
    input  io_enq_bits_lock,
    input [3:0] io_enq_bits_cache,
    input [2:0] io_enq_bits_prot,
    input [3:0] io_enq_bits_qos,
    input [3:0] io_enq_bits_region,
    input [5:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_len,
    output[2:0] io_deq_bits_size,
    output[1:0] io_deq_bits_burst,
    output io_deq_bits_lock,
    output[3:0] io_deq_bits_cache,
    output[2:0] io_deq_bits_prot,
    output[3:0] io_deq_bits_qos,
    output[3:0] io_deq_bits_region,
    output[5:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T37;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T38;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T39;
  wire T8;
  wire T9;
  wire T10;
  wire[67:0] T11;
  reg [67:0] ram [1:0];
  wire[67:0] T12;
  wire[67:0] T13;
  wire[67:0] T14;
  wire[21:0] T15;
  wire[10:0] T16;
  wire[6:0] T17;
  wire[10:0] T18;
  wire[6:0] T19;
  wire[45:0] T20;
  wire[5:0] T21;
  wire[2:0] T22;
  wire[39:0] T23;
  wire[5:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[2:0] T27;
  wire[3:0] T28;
  wire T29;
  wire[1:0] T30;
  wire[2:0] T31;
  wire[7:0] T32;
  wire[31:0] T33;
  wire T34;
  wire empty;
  wire T35;
  wire T36;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T37 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T38 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T39 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T20, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_region, T17};
  assign T17 = {io_enq_bits_id, io_enq_bits_user};
  assign T18 = {io_enq_bits_cache, T19};
  assign T19 = {io_enq_bits_prot, io_enq_bits_qos};
  assign T20 = {T23, T21};
  assign T21 = {io_enq_bits_size, T22};
  assign T22 = {io_enq_bits_burst, io_enq_bits_lock};
  assign T23 = {io_enq_bits_addr, io_enq_bits_len};
  assign io_deq_bits_id = T24;
  assign T24 = T11[3'h6:1'h1];
  assign io_deq_bits_region = T25;
  assign T25 = T11[4'ha:3'h7];
  assign io_deq_bits_qos = T26;
  assign T26 = T11[4'he:4'hb];
  assign io_deq_bits_prot = T27;
  assign T27 = T11[5'h11:4'hf];
  assign io_deq_bits_cache = T28;
  assign T28 = T11[5'h15:5'h12];
  assign io_deq_bits_lock = T29;
  assign T29 = T11[5'h16];
  assign io_deq_bits_burst = T30;
  assign T30 = T11[5'h18:5'h17];
  assign io_deq_bits_size = T31;
  assign T31 = T11[5'h1b:5'h19];
  assign io_deq_bits_len = T32;
  assign T32 = T11[6'h23:5'h1c];
  assign io_deq_bits_addr = T33;
  assign T33 = T11[7'h43:6'h24];
  assign io_deq_valid = T34;
  assign T34 = empty ^ 1'h1;
  assign empty = ptr_match & T35;
  assign T35 = maybe_full ^ 1'h1;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_19(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [5:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[5:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[5:0] T10;
  reg [5:0] ram [1:0];
  wire[5:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module NastiErrorSlave(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [5:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[5:0] io_b_bits_id,
    //output io_b_bits_user
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [5:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[5:0] io_r_bits_id
    //output io_r_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[31:0] T3;
  wire[247:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire[239:0] T9;
  wire T10;
  wire T11;
  reg  draining;
  wire T39;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg [7:0] beats_left;
  wire[7:0] T40;
  wire[7:0] T22;
  wire[7:0] T23;
  wire T24;
  wire T25;
  reg  responding;
  wire T41;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire r_queue_io_enq_ready;
  wire r_queue_io_deq_valid;
  wire[7:0] r_queue_io_deq_bits_len;
  wire[5:0] r_queue_io_deq_bits_id;
  wire b_queue_io_enq_ready;
  wire b_queue_io_deq_valid;
  wire[5:0] b_queue_io_deq_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    draining = {1{$random}};
    beats_left = {1{$random}};
    responding = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_r_bits_user = {1{$random}};
//  assign io_b_bits_user = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T2 & T1;
  assign T1 = reset ^ 1'h1;
  assign T2 = io_aw_ready & io_aw_valid;
  assign T3 = io_aw_bits_addr;
  assign T5 = T7 & T6;
  assign T6 = reset ^ 1'h1;
  assign T7 = io_ar_ready & io_ar_valid;
  assign T8 = io_ar_bits_addr;
  assign T10 = io_b_ready & T11;
  assign T11 = draining ^ 1'h1;
  assign T39 = reset ? 1'h0 : T12;
  assign T12 = T15 ? 1'h0 : T13;
  assign T13 = T14 ? 1'h1 : draining;
  assign T14 = io_aw_ready & io_aw_valid;
  assign T15 = T16 & io_w_bits_last;
  assign T16 = io_w_ready & io_w_valid;
  assign T17 = io_aw_valid & T18;
  assign T18 = draining ^ 1'h1;
  assign T19 = T20 & io_r_bits_last;
  assign T20 = io_r_ready & io_r_valid;
  assign io_r_bits_id = r_queue_io_deq_bits_id;
  assign io_r_bits_last = T21;
  assign T21 = beats_left == 8'h0;
  assign T40 = reset ? 8'h0 : T22;
  assign T22 = T32 ? T31 : T23;
  assign T23 = T24 ? r_queue_io_deq_bits_len : beats_left;
  assign T24 = T25 & r_queue_io_deq_valid;
  assign T25 = responding ^ 1'h1;
  assign T41 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h0 : T27;
  assign T27 = T24 ? 1'h1 : responding;
  assign T28 = T30 & T29;
  assign T29 = beats_left == 8'h0;
  assign T30 = io_r_ready & io_r_valid;
  assign T31 = beats_left - 8'h1;
  assign T32 = T30 & T33;
  assign T33 = T29 ^ 1'h1;
  assign io_r_bits_data = 64'h0;
  assign io_r_bits_resp = 2'h3;
  assign io_r_valid = T34;
  assign T34 = r_queue_io_deq_valid & responding;
  assign io_ar_ready = r_queue_io_enq_ready;
  assign io_b_bits_id = b_queue_io_deq_bits;
  assign io_b_bits_resp = 2'h3;
  assign io_b_valid = T35;
  assign T35 = b_queue_io_deq_valid & T36;
  assign T36 = draining ^ 1'h1;
  assign io_w_ready = draining;
  assign io_aw_ready = T37;
  assign T37 = b_queue_io_enq_ready & T38;
  assign T38 = draining ^ 1'h1;
  Queue_2 r_queue(.clk(clk), .reset(reset),
       .io_enq_ready( r_queue_io_enq_ready ),
       .io_enq_valid( io_ar_valid ),
       .io_enq_bits_addr( io_ar_bits_addr ),
       .io_enq_bits_len( io_ar_bits_len ),
       .io_enq_bits_size( io_ar_bits_size ),
       .io_enq_bits_burst( io_ar_bits_burst ),
       .io_enq_bits_lock( io_ar_bits_lock ),
       .io_enq_bits_cache( io_ar_bits_cache ),
       .io_enq_bits_prot( io_ar_bits_prot ),
       .io_enq_bits_qos( io_ar_bits_qos ),
       .io_enq_bits_region( io_ar_bits_region ),
       .io_enq_bits_id( io_ar_bits_id ),
       .io_enq_bits_user( io_ar_bits_user ),
       .io_deq_ready( T19 ),
       .io_deq_valid( r_queue_io_deq_valid ),
       //.io_deq_bits_addr(  )
       .io_deq_bits_len( r_queue_io_deq_bits_len ),
       //.io_deq_bits_size(  )
       //.io_deq_bits_burst(  )
       //.io_deq_bits_lock(  )
       //.io_deq_bits_cache(  )
       //.io_deq_bits_prot(  )
       //.io_deq_bits_qos(  )
       //.io_deq_bits_region(  )
       .io_deq_bits_id( r_queue_io_deq_bits_id )
       //.io_deq_bits_user(  )
       //.io_count(  )
  );
  Queue_19 b_queue(.clk(clk), .reset(reset),
       .io_enq_ready( b_queue_io_enq_ready ),
       .io_enq_valid( T17 ),
       .io_enq_bits( io_aw_bits_id ),
       .io_deq_ready( T10 ),
       .io_deq_valid( b_queue_io_deq_valid ),
       .io_deq_bits( b_queue_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      draining <= 1'h0;
    end else if(T15) begin
      draining <= 1'h0;
    end else if(T14) begin
      draining <= 1'h1;
    end
    if(reset) begin
      beats_left <= 8'h0;
    end else if(T32) begin
      beats_left <= T31;
    end else if(T24) begin
      beats_left <= r_queue_io_deq_bits_len;
    end
    if(reset) begin
      responding <= 1'h0;
    end else if(T28) begin
      responding <= 1'h0;
    end else if(T24) begin
      responding <= 1'h1;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T5)
        $fwrite(32'h80000002, "Invalid read address %h\n", T8);
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "Invalid write address %h\n", T3);
// synthesis translate_on
`endif
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [5:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [5:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [5:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[5:0] io_out_bits_id,
    output io_out_bits_user,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[5:0] T14;
  wire[5:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_user = T9;
  assign T9 = T13 ? io_in_2_bits_user : T10;
  assign T10 = T11 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T11 = T12[1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1];
  assign io_out_bits_id = T14;
  assign T14 = T17 ? io_in_2_bits_id : T15;
  assign T15 = T16 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T16 = T12[1'h0];
  assign T17 = T12[1'h1];
  assign io_out_bits_resp = T18;
  assign T18 = T21 ? io_in_2_bits_resp : T19;
  assign T19 = T20 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T20 = T12[1'h0];
  assign T21 = T12[1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0];
  assign T25 = T12[1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module JunctionsPeekingArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [63:0] io_in_2_bits_data,
    input  io_in_2_bits_last,
    input [5:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_last,
    input [5:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_last,
    input [5:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[63:0] io_out_bits_data,
    output io_out_bits_last,
    output[5:0] io_out_bits_id,
    output io_out_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] chosen;
  wire[1:0] choice;
  wire[1:0] T4;
  wire[1:0] T5;
  reg [1:0] T6;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  reg [1:0] T14;
  wire[1:0] T15;
  reg [1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire[1:0] T34;
  reg [1:0] T35;
  wire[1:0] T36;
  reg [1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  reg [1:0] lockIdx;
  wire[1:0] T88;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire T57;
  reg  locked;
  wire T89;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_user = T0;
  assign T0 = T61 ? io_in_2_bits_user : T1;
  assign T1 = T2 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T2 = T3[1'h0];
  assign T3 = chosen;
  assign chosen = locked ? lockIdx : choice;
  assign choice = T40 ? T34 : T4;
  assign T4 = T19 ? T13 : T5;
  assign T5 = T12 ? T10 : T6;
  always @(*) case (T8)
    0: T6 = 2'h0;
    1: T6 = 2'h1;
    2: T6 = 2'h2;
    default: begin
      T6 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T6 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T8 = T9 - 2'h1;
  assign T9 = lockIdx + 2'h1;
  always @(*) case (T11)
    0: T10 = 2'h0;
    1: T10 = 2'h1;
    2: T10 = 2'h2;
    default: begin
      T10 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T10 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T11 = 2'h2 + T9;
  assign T12 = T9 < 2'h1;
  assign T13 = T18 ? T16 : T14;
  always @(*) case (T15)
    0: T14 = 2'h0;
    1: T14 = 2'h1;
    2: T14 = 2'h2;
    default: begin
      T14 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T14 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T15 = T9 - 2'h2;
  always @(*) case (T17)
    0: T16 = 2'h0;
    1: T16 = 2'h1;
    2: T16 = 2'h2;
    default: begin
      T16 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T16 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T17 = 2'h1 + T9;
  assign T18 = T9 < 2'h2;
  assign T19 = T33 ? T27 : T20;
  assign T20 = T26 ? io_in_2_valid : T21;
  assign T21 = T22 ? io_in_1_valid : io_in_0_valid;
  assign T22 = T23[1'h0];
  assign T23 = T24;
  assign T24 = T25 - 2'h2;
  assign T25 = lockIdx + 2'h1;
  assign T26 = T23[1'h1];
  assign T27 = T32 ? io_in_2_valid : T28;
  assign T28 = T29 ? io_in_1_valid : io_in_0_valid;
  assign T29 = T30[1'h0];
  assign T30 = T31;
  assign T31 = 2'h1 + T25;
  assign T32 = T30[1'h1];
  assign T33 = T25 < 2'h2;
  assign T34 = T39 ? T37 : T35;
  always @(*) case (T36)
    0: T35 = 2'h0;
    1: T35 = 2'h1;
    2: T35 = 2'h2;
    default: begin
      T35 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T35 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T36 = T9 - 2'h3;
  always @(*) case (T38)
    0: T37 = 2'h0;
    1: T37 = 2'h1;
    2: T37 = 2'h2;
    default: begin
      T37 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T37 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T38 = 2'h0 + T9;
  assign T39 = T9 < 2'h3;
  assign T40 = T53 ? T47 : T41;
  assign T41 = T46 ? io_in_2_valid : T42;
  assign T42 = T43 ? io_in_1_valid : io_in_0_valid;
  assign T43 = T44[1'h0];
  assign T44 = T45;
  assign T45 = T25 - 2'h3;
  assign T46 = T44[1'h1];
  assign T47 = T52 ? io_in_2_valid : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T50[1'h0];
  assign T50 = T51;
  assign T51 = 2'h0 + T25;
  assign T52 = T50[1'h1];
  assign T53 = T25 < 2'h3;
  assign T88 = reset ? 2'h0 : T54;
  assign T54 = T55 ? choice : lockIdx;
  assign T55 = T57 & T56;
  assign T56 = locked ^ 1'h1;
  assign T57 = io_out_ready & io_out_valid;
  assign T89 = reset ? 1'h0 : T58;
  assign T58 = T60 ? 1'h0 : T59;
  assign T59 = T55 ? 1'h1 : locked;
  assign T60 = T57 & io_out_bits_last;
  assign T61 = T3[1'h1];
  assign io_out_bits_id = T62;
  assign T62 = T65 ? io_in_2_bits_id : T63;
  assign T63 = T64 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T64 = T3[1'h0];
  assign T65 = T3[1'h1];
  assign io_out_bits_last = T66;
  assign T66 = T69 ? io_in_2_bits_last : T67;
  assign T67 = T68 ? io_in_1_bits_last : io_in_0_bits_last;
  assign T68 = T3[1'h0];
  assign T69 = T3[1'h1];
  assign io_out_bits_data = T70;
  assign T70 = T73 ? io_in_2_bits_data : T71;
  assign T71 = T72 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T72 = T3[1'h0];
  assign T73 = T3[1'h1];
  assign io_out_bits_resp = T74;
  assign T74 = T77 ? io_in_2_bits_resp : T75;
  assign T75 = T76 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T76 = T3[1'h0];
  assign T77 = T3[1'h1];
  assign io_out_valid = T78;
  assign T78 = T81 ? io_in_2_valid : T79;
  assign T79 = T80 ? io_in_1_valid : io_in_0_valid;
  assign T80 = T3[1'h0];
  assign T81 = T3[1'h1];
  assign io_in_0_ready = T82;
  assign T82 = io_out_ready & T83;
  assign T83 = chosen == 2'h0;
  assign io_in_1_ready = T84;
  assign T84 = io_out_ready & T85;
  assign T85 = chosen == 2'h1;
  assign io_in_2_ready = T86;
  assign T86 = io_out_ready & T87;
  assign T87 = chosen == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h0;
    end else if(T55) begin
      lockIdx <= choice;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T60) begin
      locked <= 1'h0;
    end else if(T55) begin
      locked <= 1'h1;
    end
  end
endmodule

module NastiRouter_0(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [5:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[5:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [5:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[5:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[5:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [5:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[5:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [5:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[5:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [5:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[5:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [5:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[1:0] ar_route;
  wire[1:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[32:0] T55;
  wire T8;
  wire T9;
  wire w_invalid;
  wire T10;
  wire[1:0] aw_route;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[32:0] T56;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  R21;
  wire T57;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  R32;
  wire T58;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire ar_ready;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire w_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire aw_ready;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[5:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[5:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[5:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[5:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R21 = {1{$random}};
    R32 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 2'h0;
  assign ar_route = T2;
  assign T2 = {T6, T3};
  assign T3 = T5 & T4;
  assign T4 = io_master_ar_bits_addr < 32'h80000000;
  assign T5 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T6 = T8 & T7;
  assign T7 = T55 < 33'h100000000;
  assign T55 = {1'h0, io_master_ar_bits_addr};
  assign T8 = 32'h80000000 <= io_master_ar_bits_addr;
  assign T9 = w_invalid & io_master_aw_valid;
  assign w_invalid = T10 ^ 1'h1;
  assign T10 = aw_route != 2'h0;
  assign aw_route = T11;
  assign T11 = {T15, T12};
  assign T12 = T14 & T13;
  assign T13 = io_master_aw_bits_addr < 32'h80000000;
  assign T14 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T15 = T17 & T16;
  assign T16 = T56 < 33'h100000000;
  assign T56 = {1'h0, io_master_aw_bits_addr};
  assign T17 = 32'h80000000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T18;
  assign T18 = io_master_ar_valid & T19;
  assign T19 = ar_route[1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T20;
  assign T20 = io_master_w_valid & R21;
  assign T57 = reset ? 1'h0 : T22;
  assign T22 = T25 ? 1'h0 : T23;
  assign T23 = T24 ? 1'h1 : R21;
  assign T24 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T25 = T26 & io_slave_0_w_bits_last;
  assign T26 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T27;
  assign T27 = io_master_aw_valid & T28;
  assign T28 = aw_route[1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T29;
  assign T29 = io_master_ar_valid & T30;
  assign T30 = ar_route[1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T31;
  assign T31 = io_master_w_valid & R32;
  assign T58 = reset ? 1'h0 : T33;
  assign T33 = T36 ? 1'h0 : T34;
  assign T34 = T35 ? 1'h1 : R32;
  assign T35 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T36 = T37 & io_slave_1_w_bits_last;
  assign T37 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T38;
  assign T38 = io_master_aw_valid & T39;
  assign T39 = aw_route[1'h1];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T40;
  assign T40 = ar_ready | T41;
  assign T41 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T44 | T42;
  assign T42 = io_slave_1_ar_ready & T43;
  assign T43 = ar_route[1'h1];
  assign T44 = io_slave_0_ar_ready & T45;
  assign T45 = ar_route[1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T46;
  assign T46 = w_ready | err_slave_io_w_ready;
  assign w_ready = T48 | T47;
  assign T47 = io_slave_1_w_ready & R32;
  assign T48 = io_slave_0_w_ready & R21;
  assign io_master_aw_ready = T49;
  assign T49 = aw_ready | T50;
  assign T50 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T53 | T51;
  assign T51 = io_slave_1_aw_ready & T52;
  assign T52 = aw_route[1'h1];
  assign T53 = io_slave_0_aw_ready & T54;
  assign T54 = aw_route[1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T9 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_2_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_2_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_4 b_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( err_slave_io_b_valid ),
       .io_in_2_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_2_bits_id( err_slave_io_b_bits_id ),
       //.io_in_2_bits_user(  )
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_2_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter_0 r_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( err_slave_io_r_valid ),
       .io_in_2_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_2_bits_data( err_slave_io_r_bits_data ),
       .io_in_2_bits_last( err_slave_io_r_bits_last ),
       .io_in_2_bits_id( err_slave_io_r_bits_id ),
       //.io_in_2_bits_user(  )
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_2_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R21 <= 1'h0;
    end else if(T25) begin
      R21 <= 1'h0;
    end else if(T24) begin
      R21 <= 1'h1;
    end
    if(reset) begin
      R32 <= 1'h0;
    end else if(T36) begin
      R32 <= 1'h0;
    end else if(T35) begin
      R32 <= 1'h1;
    end
  end
endmodule

module RRArbiter_5(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_addr,
    input [7:0] io_in_1_bits_len,
    input [2:0] io_in_1_bits_size,
    input [1:0] io_in_1_bits_burst,
    input  io_in_1_bits_lock,
    input [3:0] io_in_1_bits_cache,
    input [2:0] io_in_1_bits_prot,
    input [3:0] io_in_1_bits_qos,
    input [3:0] io_in_1_bits_region,
    input [5:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_len,
    input [2:0] io_in_0_bits_size,
    input [1:0] io_in_0_bits_burst,
    input  io_in_0_bits_lock,
    input [3:0] io_in_0_bits_cache,
    input [2:0] io_in_0_bits_prot,
    input [3:0] io_in_0_bits_qos,
    input [3:0] io_in_0_bits_region,
    input [5:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_addr,
    output[7:0] io_out_bits_len,
    output[2:0] io_out_bits_size,
    output[1:0] io_out_bits_burst,
    output io_out_bits_lock,
    output[3:0] io_out_bits_cache,
    output[2:0] io_out_bits_prot,
    output[3:0] io_out_bits_qos,
    output[3:0] io_out_bits_region,
    output[5:0] io_out_bits_id,
    output io_out_bits_user,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T35;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[5:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[2:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire[2:0] T14;
  wire[7:0] T15;
  wire[31:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T35 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_user = T5;
  assign T5 = T6 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T6 = chosen;
  assign io_out_bits_id = T7;
  assign T7 = T6 ? io_in_1_bits_id : io_in_0_bits_id;
  assign io_out_bits_region = T8;
  assign T8 = T6 ? io_in_1_bits_region : io_in_0_bits_region;
  assign io_out_bits_qos = T9;
  assign T9 = T6 ? io_in_1_bits_qos : io_in_0_bits_qos;
  assign io_out_bits_prot = T10;
  assign T10 = T6 ? io_in_1_bits_prot : io_in_0_bits_prot;
  assign io_out_bits_cache = T11;
  assign T11 = T6 ? io_in_1_bits_cache : io_in_0_bits_cache;
  assign io_out_bits_lock = T12;
  assign T12 = T6 ? io_in_1_bits_lock : io_in_0_bits_lock;
  assign io_out_bits_burst = T13;
  assign T13 = T6 ? io_in_1_bits_burst : io_in_0_bits_burst;
  assign io_out_bits_size = T14;
  assign T14 = T6 ? io_in_1_bits_size : io_in_0_bits_size;
  assign io_out_bits_len = T15;
  assign T15 = T6 ? io_in_1_bits_len : io_in_0_bits_len;
  assign io_out_bits_addr = T16;
  assign T16 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T17;
  assign T17 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T18;
  assign T18 = T19 & io_out_ready;
  assign T19 = T26 | T20;
  assign T20 = T21 ^ 1'h1;
  assign T21 = T24 | T22;
  assign T22 = io_in_1_valid & T23;
  assign T23 = last_grant < 1'h1;
  assign T24 = io_in_0_valid & T25;
  assign T25 = last_grant < 1'h0;
  assign T26 = last_grant < 1'h0;
  assign io_in_1_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T32 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_0_valid;
  assign T31 = T24 | T22;
  assign T32 = T34 & T33;
  assign T33 = last_grant < 1'h1;
  assign T34 = T24 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module NastiArbiter_1(input clk, input reset,
    output io_master_1_aw_ready,
    input  io_master_1_aw_valid,
    input [31:0] io_master_1_aw_bits_addr,
    input [7:0] io_master_1_aw_bits_len,
    input [2:0] io_master_1_aw_bits_size,
    input [1:0] io_master_1_aw_bits_burst,
    input  io_master_1_aw_bits_lock,
    input [3:0] io_master_1_aw_bits_cache,
    input [2:0] io_master_1_aw_bits_prot,
    input [3:0] io_master_1_aw_bits_qos,
    input [3:0] io_master_1_aw_bits_region,
    input [5:0] io_master_1_aw_bits_id,
    input  io_master_1_aw_bits_user,
    output io_master_1_w_ready,
    input  io_master_1_w_valid,
    input [63:0] io_master_1_w_bits_data,
    input  io_master_1_w_bits_last,
    input [7:0] io_master_1_w_bits_strb,
    input  io_master_1_w_bits_user,
    input  io_master_1_b_ready,
    output io_master_1_b_valid,
    output[1:0] io_master_1_b_bits_resp,
    output[5:0] io_master_1_b_bits_id,
    output io_master_1_b_bits_user,
    output io_master_1_ar_ready,
    input  io_master_1_ar_valid,
    input [31:0] io_master_1_ar_bits_addr,
    input [7:0] io_master_1_ar_bits_len,
    input [2:0] io_master_1_ar_bits_size,
    input [1:0] io_master_1_ar_bits_burst,
    input  io_master_1_ar_bits_lock,
    input [3:0] io_master_1_ar_bits_cache,
    input [2:0] io_master_1_ar_bits_prot,
    input [3:0] io_master_1_ar_bits_qos,
    input [3:0] io_master_1_ar_bits_region,
    input [5:0] io_master_1_ar_bits_id,
    input  io_master_1_ar_bits_user,
    input  io_master_1_r_ready,
    output io_master_1_r_valid,
    output[1:0] io_master_1_r_bits_resp,
    output[63:0] io_master_1_r_bits_data,
    output io_master_1_r_bits_last,
    output[5:0] io_master_1_r_bits_id,
    output io_master_1_r_bits_user,
    output io_master_0_aw_ready,
    input  io_master_0_aw_valid,
    input [31:0] io_master_0_aw_bits_addr,
    input [7:0] io_master_0_aw_bits_len,
    input [2:0] io_master_0_aw_bits_size,
    input [1:0] io_master_0_aw_bits_burst,
    input  io_master_0_aw_bits_lock,
    input [3:0] io_master_0_aw_bits_cache,
    input [2:0] io_master_0_aw_bits_prot,
    input [3:0] io_master_0_aw_bits_qos,
    input [3:0] io_master_0_aw_bits_region,
    input [5:0] io_master_0_aw_bits_id,
    input  io_master_0_aw_bits_user,
    output io_master_0_w_ready,
    input  io_master_0_w_valid,
    input [63:0] io_master_0_w_bits_data,
    input  io_master_0_w_bits_last,
    input [7:0] io_master_0_w_bits_strb,
    input  io_master_0_w_bits_user,
    input  io_master_0_b_ready,
    output io_master_0_b_valid,
    output[1:0] io_master_0_b_bits_resp,
    output[5:0] io_master_0_b_bits_id,
    output io_master_0_b_bits_user,
    output io_master_0_ar_ready,
    input  io_master_0_ar_valid,
    input [31:0] io_master_0_ar_bits_addr,
    input [7:0] io_master_0_ar_bits_len,
    input [2:0] io_master_0_ar_bits_size,
    input [1:0] io_master_0_ar_bits_burst,
    input  io_master_0_ar_bits_lock,
    input [3:0] io_master_0_ar_bits_cache,
    input [2:0] io_master_0_ar_bits_prot,
    input [3:0] io_master_0_ar_bits_qos,
    input [3:0] io_master_0_ar_bits_region,
    input [5:0] io_master_0_ar_bits_id,
    input  io_master_0_ar_bits_user,
    input  io_master_0_r_ready,
    output io_master_0_r_valid,
    output[1:0] io_master_0_r_bits_resp,
    output[63:0] io_master_0_r_bits_data,
    output io_master_0_r_bits_last,
    output[5:0] io_master_0_r_bits_id,
    output io_master_0_r_bits_user,
    input  io_slave_aw_ready,
    output io_slave_aw_valid,
    output[31:0] io_slave_aw_bits_addr,
    output[7:0] io_slave_aw_bits_len,
    output[2:0] io_slave_aw_bits_size,
    output[1:0] io_slave_aw_bits_burst,
    output io_slave_aw_bits_lock,
    output[3:0] io_slave_aw_bits_cache,
    output[2:0] io_slave_aw_bits_prot,
    output[3:0] io_slave_aw_bits_qos,
    output[3:0] io_slave_aw_bits_region,
    output[5:0] io_slave_aw_bits_id,
    output io_slave_aw_bits_user,
    input  io_slave_w_ready,
    output io_slave_w_valid,
    output[63:0] io_slave_w_bits_data,
    output io_slave_w_bits_last,
    output[7:0] io_slave_w_bits_strb,
    output io_slave_w_bits_user,
    output io_slave_b_ready,
    input  io_slave_b_valid,
    input [1:0] io_slave_b_bits_resp,
    input [5:0] io_slave_b_bits_id,
    input  io_slave_b_bits_user,
    input  io_slave_ar_ready,
    output io_slave_ar_valid,
    output[31:0] io_slave_ar_bits_addr,
    output[7:0] io_slave_ar_bits_len,
    output[2:0] io_slave_ar_bits_size,
    output[1:0] io_slave_ar_bits_burst,
    output io_slave_ar_bits_lock,
    output[3:0] io_slave_ar_bits_cache,
    output[2:0] io_slave_ar_bits_prot,
    output[3:0] io_slave_ar_bits_qos,
    output[3:0] io_slave_ar_bits_region,
    output[5:0] io_slave_ar_bits_id,
    output io_slave_ar_bits_user,
    output io_slave_r_ready,
    input  io_slave_r_valid,
    input [1:0] io_slave_r_bits_resp,
    input [63:0] io_slave_r_bits_data,
    input  io_slave_r_bits_last,
    input [5:0] io_slave_r_bits_id,
    input  io_slave_r_bits_user
);

  wire T0;
  reg  R1;
  wire T48;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[5:0] T49;
  wire[6:0] T7;
  wire[5:0] T50;
  wire[6:0] T8;
  wire[5:0] T51;
  wire[6:0] T9;
  wire[5:0] T52;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg  R19;
  wire T20;
  wire[7:0] T21;
  wire T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[5:0] T53;
  wire[4:0] T28;
  wire T29;
  wire T30;
  wire[5:0] T54;
  wire[4:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[5:0] T55;
  wire[4:0] T38;
  wire T39;
  wire T40;
  wire[5:0] T56;
  wire[4:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[31:0] RRArbiter_io_out_bits_addr;
  wire[7:0] RRArbiter_io_out_bits_len;
  wire[2:0] RRArbiter_io_out_bits_size;
  wire[1:0] RRArbiter_io_out_bits_burst;
  wire RRArbiter_io_out_bits_lock;
  wire[3:0] RRArbiter_io_out_bits_cache;
  wire[2:0] RRArbiter_io_out_bits_prot;
  wire[3:0] RRArbiter_io_out_bits_qos;
  wire[3:0] RRArbiter_io_out_bits_region;
  wire[5:0] RRArbiter_io_out_bits_id;
  wire RRArbiter_io_out_bits_user;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[31:0] RRArbiter_1_io_out_bits_addr;
  wire[7:0] RRArbiter_1_io_out_bits_len;
  wire[2:0] RRArbiter_1_io_out_bits_size;
  wire[1:0] RRArbiter_1_io_out_bits_burst;
  wire RRArbiter_1_io_out_bits_lock;
  wire[3:0] RRArbiter_1_io_out_bits_cache;
  wire[2:0] RRArbiter_1_io_out_bits_prot;
  wire[3:0] RRArbiter_1_io_out_bits_qos;
  wire[3:0] RRArbiter_1_io_out_bits_region;
  wire[5:0] RRArbiter_1_io_out_bits_id;
  wire RRArbiter_1_io_out_bits_user;
  wire RRArbiter_1_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R19 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_slave_aw_ready & R1;
  assign T48 = reset ? 1'h1 : T2;
  assign T2 = T5 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : R1;
  assign T4 = T0 & RRArbiter_1_io_out_valid;
  assign T5 = T6 & io_slave_w_bits_last;
  assign T6 = io_slave_w_ready & io_slave_w_valid;
  assign T49 = T7[3'h5:1'h0];
  assign T7 = {io_master_0_aw_bits_id, 1'h0};
  assign T50 = T8[3'h5:1'h0];
  assign T8 = {io_master_1_aw_bits_id, 1'h1};
  assign T51 = T9[3'h5:1'h0];
  assign T9 = {io_master_0_ar_bits_id, 1'h0};
  assign T52 = T10[3'h5:1'h0];
  assign T10 = {io_master_1_ar_bits_id, 1'h1};
  assign io_slave_r_ready = T11;
  assign T11 = T12 ? io_master_1_r_ready : io_master_0_r_ready;
  assign T12 = T13;
  assign T13 = io_slave_r_bits_id[1'h0];
  assign io_slave_ar_bits_user = RRArbiter_io_out_bits_user;
  assign io_slave_ar_bits_id = RRArbiter_io_out_bits_id;
  assign io_slave_ar_bits_region = RRArbiter_io_out_bits_region;
  assign io_slave_ar_bits_qos = RRArbiter_io_out_bits_qos;
  assign io_slave_ar_bits_prot = RRArbiter_io_out_bits_prot;
  assign io_slave_ar_bits_cache = RRArbiter_io_out_bits_cache;
  assign io_slave_ar_bits_lock = RRArbiter_io_out_bits_lock;
  assign io_slave_ar_bits_burst = RRArbiter_io_out_bits_burst;
  assign io_slave_ar_bits_size = RRArbiter_io_out_bits_size;
  assign io_slave_ar_bits_len = RRArbiter_io_out_bits_len;
  assign io_slave_ar_bits_addr = RRArbiter_io_out_bits_addr;
  assign io_slave_ar_valid = RRArbiter_io_out_valid;
  assign io_slave_b_ready = T14;
  assign T14 = T15 ? io_master_1_b_ready : io_master_0_b_ready;
  assign T15 = T16;
  assign T16 = io_slave_b_bits_id[1'h0];
  assign io_slave_w_bits_user = T17;
  assign T17 = T18 ? io_master_1_w_bits_user : io_master_0_w_bits_user;
  assign T18 = R19;
  assign T20 = T4 ? RRArbiter_1_io_chosen : R19;
  assign io_slave_w_bits_strb = T21;
  assign T21 = T18 ? io_master_1_w_bits_strb : io_master_0_w_bits_strb;
  assign io_slave_w_bits_last = T22;
  assign T22 = T18 ? io_master_1_w_bits_last : io_master_0_w_bits_last;
  assign io_slave_w_bits_data = T23;
  assign T23 = T18 ? io_master_1_w_bits_data : io_master_0_w_bits_data;
  assign io_slave_w_valid = T24;
  assign T24 = T26 & T25;
  assign T25 = R1 ^ 1'h1;
  assign T26 = T18 ? io_master_1_w_valid : io_master_0_w_valid;
  assign io_slave_aw_bits_user = RRArbiter_1_io_out_bits_user;
  assign io_slave_aw_bits_id = RRArbiter_1_io_out_bits_id;
  assign io_slave_aw_bits_region = RRArbiter_1_io_out_bits_region;
  assign io_slave_aw_bits_qos = RRArbiter_1_io_out_bits_qos;
  assign io_slave_aw_bits_prot = RRArbiter_1_io_out_bits_prot;
  assign io_slave_aw_bits_cache = RRArbiter_1_io_out_bits_cache;
  assign io_slave_aw_bits_lock = RRArbiter_1_io_out_bits_lock;
  assign io_slave_aw_bits_burst = RRArbiter_1_io_out_bits_burst;
  assign io_slave_aw_bits_size = RRArbiter_1_io_out_bits_size;
  assign io_slave_aw_bits_len = RRArbiter_1_io_out_bits_len;
  assign io_slave_aw_bits_addr = RRArbiter_1_io_out_bits_addr;
  assign io_slave_aw_valid = T27;
  assign T27 = RRArbiter_1_io_out_valid & R1;
  assign io_master_0_r_bits_user = io_slave_r_bits_user;
  assign io_master_0_r_bits_id = T53;
  assign T53 = {1'h0, T28};
  assign T28 = io_slave_r_bits_id >> 1'h1;
  assign io_master_0_r_bits_last = io_slave_r_bits_last;
  assign io_master_0_r_bits_data = io_slave_r_bits_data;
  assign io_master_0_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_0_r_valid = T29;
  assign T29 = io_slave_r_valid & T30;
  assign T30 = T13 == 1'h0;
  assign io_master_0_ar_ready = RRArbiter_io_in_0_ready;
  assign io_master_0_b_bits_user = io_slave_b_bits_user;
  assign io_master_0_b_bits_id = T54;
  assign T54 = {1'h0, T31};
  assign T31 = io_slave_b_bits_id >> 1'h1;
  assign io_master_0_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_0_b_valid = T32;
  assign T32 = io_slave_b_valid & T33;
  assign T33 = T16 == 1'h0;
  assign io_master_0_w_ready = T34;
  assign T34 = T36 & T35;
  assign T35 = R1 ^ 1'h1;
  assign T36 = io_slave_w_ready & T37;
  assign T37 = R19 == 1'h0;
  assign io_master_0_aw_ready = RRArbiter_1_io_in_0_ready;
  assign io_master_1_r_bits_user = io_slave_r_bits_user;
  assign io_master_1_r_bits_id = T55;
  assign T55 = {1'h0, T38};
  assign T38 = io_slave_r_bits_id >> 1'h1;
  assign io_master_1_r_bits_last = io_slave_r_bits_last;
  assign io_master_1_r_bits_data = io_slave_r_bits_data;
  assign io_master_1_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_1_r_valid = T39;
  assign T39 = io_slave_r_valid & T40;
  assign T40 = T13 == 1'h1;
  assign io_master_1_ar_ready = RRArbiter_io_in_1_ready;
  assign io_master_1_b_bits_user = io_slave_b_bits_user;
  assign io_master_1_b_bits_id = T56;
  assign T56 = {1'h0, T41};
  assign T41 = io_slave_b_bits_id >> 1'h1;
  assign io_master_1_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_1_b_valid = T42;
  assign T42 = io_slave_b_valid & T43;
  assign T43 = T16 == 1'h1;
  assign io_master_1_w_ready = T44;
  assign T44 = T46 & T45;
  assign T45 = R1 ^ 1'h1;
  assign T46 = io_slave_w_ready & T47;
  assign T47 = R19 == 1'h1;
  assign io_master_1_aw_ready = RRArbiter_1_io_in_1_ready;
  RRArbiter_5 RRArbiter(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_master_1_ar_valid ),
       .io_in_1_bits_addr( io_master_1_ar_bits_addr ),
       .io_in_1_bits_len( io_master_1_ar_bits_len ),
       .io_in_1_bits_size( io_master_1_ar_bits_size ),
       .io_in_1_bits_burst( io_master_1_ar_bits_burst ),
       .io_in_1_bits_lock( io_master_1_ar_bits_lock ),
       .io_in_1_bits_cache( io_master_1_ar_bits_cache ),
       .io_in_1_bits_prot( io_master_1_ar_bits_prot ),
       .io_in_1_bits_qos( io_master_1_ar_bits_qos ),
       .io_in_1_bits_region( io_master_1_ar_bits_region ),
       .io_in_1_bits_id( T52 ),
       .io_in_1_bits_user( io_master_1_ar_bits_user ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_master_0_ar_valid ),
       .io_in_0_bits_addr( io_master_0_ar_bits_addr ),
       .io_in_0_bits_len( io_master_0_ar_bits_len ),
       .io_in_0_bits_size( io_master_0_ar_bits_size ),
       .io_in_0_bits_burst( io_master_0_ar_bits_burst ),
       .io_in_0_bits_lock( io_master_0_ar_bits_lock ),
       .io_in_0_bits_cache( io_master_0_ar_bits_cache ),
       .io_in_0_bits_prot( io_master_0_ar_bits_prot ),
       .io_in_0_bits_qos( io_master_0_ar_bits_qos ),
       .io_in_0_bits_region( io_master_0_ar_bits_region ),
       .io_in_0_bits_id( T51 ),
       .io_in_0_bits_user( io_master_0_ar_bits_user ),
       .io_out_ready( io_slave_ar_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_addr( RRArbiter_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_io_out_bits_user )
       //.io_chosen(  )
  );
  RRArbiter_5 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_master_1_aw_valid ),
       .io_in_1_bits_addr( io_master_1_aw_bits_addr ),
       .io_in_1_bits_len( io_master_1_aw_bits_len ),
       .io_in_1_bits_size( io_master_1_aw_bits_size ),
       .io_in_1_bits_burst( io_master_1_aw_bits_burst ),
       .io_in_1_bits_lock( io_master_1_aw_bits_lock ),
       .io_in_1_bits_cache( io_master_1_aw_bits_cache ),
       .io_in_1_bits_prot( io_master_1_aw_bits_prot ),
       .io_in_1_bits_qos( io_master_1_aw_bits_qos ),
       .io_in_1_bits_region( io_master_1_aw_bits_region ),
       .io_in_1_bits_id( T50 ),
       .io_in_1_bits_user( io_master_1_aw_bits_user ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_master_0_aw_valid ),
       .io_in_0_bits_addr( io_master_0_aw_bits_addr ),
       .io_in_0_bits_len( io_master_0_aw_bits_len ),
       .io_in_0_bits_size( io_master_0_aw_bits_size ),
       .io_in_0_bits_burst( io_master_0_aw_bits_burst ),
       .io_in_0_bits_lock( io_master_0_aw_bits_lock ),
       .io_in_0_bits_cache( io_master_0_aw_bits_cache ),
       .io_in_0_bits_prot( io_master_0_aw_bits_prot ),
       .io_in_0_bits_qos( io_master_0_aw_bits_qos ),
       .io_in_0_bits_region( io_master_0_aw_bits_region ),
       .io_in_0_bits_id( T49 ),
       .io_in_0_bits_user( io_master_0_aw_bits_user ),
       .io_out_ready( T0 ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_addr( RRArbiter_1_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_1_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_1_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_1_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_1_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_1_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_1_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_1_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_1_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_1_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_1_io_out_bits_user ),
       .io_chosen( RRArbiter_1_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h1;
    end else if(T5) begin
      R1 <= 1'h1;
    end else if(T4) begin
      R1 <= 1'h0;
    end
    if(T4) begin
      R19 <= RRArbiter_1_io_chosen;
    end
  end
endmodule

module NastiCrossbar_0(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [5:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[5:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [5:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[5:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [5:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[5:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [5:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[5:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[5:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [5:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[5:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [5:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[5:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [5:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[5:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [5:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiArbiter_io_master_1_aw_ready;
  wire NastiArbiter_io_master_1_w_ready;
  wire NastiArbiter_io_master_1_b_valid;
  wire[1:0] NastiArbiter_io_master_1_b_bits_resp;
  wire[5:0] NastiArbiter_io_master_1_b_bits_id;
  wire NastiArbiter_io_master_1_b_bits_user;
  wire NastiArbiter_io_master_1_ar_ready;
  wire NastiArbiter_io_master_1_r_valid;
  wire[1:0] NastiArbiter_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_1_r_bits_data;
  wire NastiArbiter_io_master_1_r_bits_last;
  wire[5:0] NastiArbiter_io_master_1_r_bits_id;
  wire NastiArbiter_io_master_1_r_bits_user;
  wire NastiArbiter_io_master_0_aw_ready;
  wire NastiArbiter_io_master_0_w_ready;
  wire NastiArbiter_io_master_0_b_valid;
  wire[1:0] NastiArbiter_io_master_0_b_bits_resp;
  wire[5:0] NastiArbiter_io_master_0_b_bits_id;
  wire NastiArbiter_io_master_0_b_bits_user;
  wire NastiArbiter_io_master_0_ar_ready;
  wire NastiArbiter_io_master_0_r_valid;
  wire[1:0] NastiArbiter_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_0_r_bits_data;
  wire NastiArbiter_io_master_0_r_bits_last;
  wire[5:0] NastiArbiter_io_master_0_r_bits_id;
  wire NastiArbiter_io_master_0_r_bits_user;
  wire NastiArbiter_io_slave_aw_valid;
  wire[31:0] NastiArbiter_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_io_slave_aw_bits_burst;
  wire NastiArbiter_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_io_slave_aw_bits_region;
  wire[5:0] NastiArbiter_io_slave_aw_bits_id;
  wire NastiArbiter_io_slave_aw_bits_user;
  wire NastiArbiter_io_slave_w_valid;
  wire[63:0] NastiArbiter_io_slave_w_bits_data;
  wire NastiArbiter_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_io_slave_w_bits_strb;
  wire NastiArbiter_io_slave_w_bits_user;
  wire NastiArbiter_io_slave_b_ready;
  wire NastiArbiter_io_slave_ar_valid;
  wire[31:0] NastiArbiter_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_io_slave_ar_bits_burst;
  wire NastiArbiter_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_io_slave_ar_bits_region;
  wire[5:0] NastiArbiter_io_slave_ar_bits_id;
  wire NastiArbiter_io_slave_ar_bits_user;
  wire NastiArbiter_io_slave_r_ready;
  wire NastiArbiter_1_io_master_1_aw_ready;
  wire NastiArbiter_1_io_master_1_w_ready;
  wire NastiArbiter_1_io_master_1_b_valid;
  wire[1:0] NastiArbiter_1_io_master_1_b_bits_resp;
  wire[5:0] NastiArbiter_1_io_master_1_b_bits_id;
  wire NastiArbiter_1_io_master_1_b_bits_user;
  wire NastiArbiter_1_io_master_1_ar_ready;
  wire NastiArbiter_1_io_master_1_r_valid;
  wire[1:0] NastiArbiter_1_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_1_r_bits_data;
  wire NastiArbiter_1_io_master_1_r_bits_last;
  wire[5:0] NastiArbiter_1_io_master_1_r_bits_id;
  wire NastiArbiter_1_io_master_1_r_bits_user;
  wire NastiArbiter_1_io_master_0_aw_ready;
  wire NastiArbiter_1_io_master_0_w_ready;
  wire NastiArbiter_1_io_master_0_b_valid;
  wire[1:0] NastiArbiter_1_io_master_0_b_bits_resp;
  wire[5:0] NastiArbiter_1_io_master_0_b_bits_id;
  wire NastiArbiter_1_io_master_0_b_bits_user;
  wire NastiArbiter_1_io_master_0_ar_ready;
  wire NastiArbiter_1_io_master_0_r_valid;
  wire[1:0] NastiArbiter_1_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_0_r_bits_data;
  wire NastiArbiter_1_io_master_0_r_bits_last;
  wire[5:0] NastiArbiter_1_io_master_0_r_bits_id;
  wire NastiArbiter_1_io_master_0_r_bits_user;
  wire NastiArbiter_1_io_slave_aw_valid;
  wire[31:0] NastiArbiter_1_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_aw_bits_burst;
  wire NastiArbiter_1_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_region;
  wire[5:0] NastiArbiter_1_io_slave_aw_bits_id;
  wire NastiArbiter_1_io_slave_aw_bits_user;
  wire NastiArbiter_1_io_slave_w_valid;
  wire[63:0] NastiArbiter_1_io_slave_w_bits_data;
  wire NastiArbiter_1_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_1_io_slave_w_bits_strb;
  wire NastiArbiter_1_io_slave_w_bits_user;
  wire NastiArbiter_1_io_slave_b_ready;
  wire NastiArbiter_1_io_slave_ar_valid;
  wire[31:0] NastiArbiter_1_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_ar_bits_burst;
  wire NastiArbiter_1_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_region;
  wire[5:0] NastiArbiter_1_io_slave_ar_bits_id;
  wire NastiArbiter_1_io_slave_ar_bits_user;
  wire NastiArbiter_1_io_slave_r_ready;
  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[5:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[5:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[5:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[5:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[5:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[5:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;
  wire NastiRouter_1_io_master_aw_ready;
  wire NastiRouter_1_io_master_w_ready;
  wire NastiRouter_1_io_master_b_valid;
  wire[1:0] NastiRouter_1_io_master_b_bits_resp;
  wire[5:0] NastiRouter_1_io_master_b_bits_id;
  wire NastiRouter_1_io_master_b_bits_user;
  wire NastiRouter_1_io_master_ar_ready;
  wire NastiRouter_1_io_master_r_valid;
  wire[1:0] NastiRouter_1_io_master_r_bits_resp;
  wire[63:0] NastiRouter_1_io_master_r_bits_data;
  wire NastiRouter_1_io_master_r_bits_last;
  wire[5:0] NastiRouter_1_io_master_r_bits_id;
  wire NastiRouter_1_io_master_r_bits_user;
  wire NastiRouter_1_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_aw_bits_burst;
  wire NastiRouter_1_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_region;
  wire[5:0] NastiRouter_1_io_slave_1_aw_bits_id;
  wire NastiRouter_1_io_slave_1_aw_bits_user;
  wire NastiRouter_1_io_slave_1_w_valid;
  wire[63:0] NastiRouter_1_io_slave_1_w_bits_data;
  wire NastiRouter_1_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_1_w_bits_strb;
  wire NastiRouter_1_io_slave_1_w_bits_user;
  wire NastiRouter_1_io_slave_1_b_ready;
  wire NastiRouter_1_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_ar_bits_burst;
  wire NastiRouter_1_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_region;
  wire[5:0] NastiRouter_1_io_slave_1_ar_bits_id;
  wire NastiRouter_1_io_slave_1_ar_bits_user;
  wire NastiRouter_1_io_slave_1_r_ready;
  wire NastiRouter_1_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_aw_bits_burst;
  wire NastiRouter_1_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_region;
  wire[5:0] NastiRouter_1_io_slave_0_aw_bits_id;
  wire NastiRouter_1_io_slave_0_aw_bits_user;
  wire NastiRouter_1_io_slave_0_w_valid;
  wire[63:0] NastiRouter_1_io_slave_0_w_bits_data;
  wire NastiRouter_1_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_0_w_bits_strb;
  wire NastiRouter_1_io_slave_0_w_bits_user;
  wire NastiRouter_1_io_slave_0_b_ready;
  wire NastiRouter_1_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_ar_bits_burst;
  wire NastiRouter_1_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_region;
  wire[5:0] NastiRouter_1_io_slave_0_ar_bits_id;
  wire NastiRouter_1_io_slave_0_ar_bits_user;
  wire NastiRouter_1_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiArbiter_io_slave_r_ready;
  assign io_slaves_0_ar_bits_user = NastiArbiter_io_slave_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiArbiter_io_slave_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiArbiter_io_slave_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiArbiter_io_slave_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiArbiter_io_slave_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiArbiter_io_slave_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiArbiter_io_slave_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiArbiter_io_slave_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiArbiter_io_slave_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiArbiter_io_slave_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiArbiter_io_slave_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiArbiter_io_slave_ar_valid;
  assign io_slaves_0_b_ready = NastiArbiter_io_slave_b_ready;
  assign io_slaves_0_w_bits_user = NastiArbiter_io_slave_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiArbiter_io_slave_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiArbiter_io_slave_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiArbiter_io_slave_w_bits_data;
  assign io_slaves_0_w_valid = NastiArbiter_io_slave_w_valid;
  assign io_slaves_0_aw_bits_user = NastiArbiter_io_slave_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiArbiter_io_slave_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiArbiter_io_slave_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiArbiter_io_slave_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiArbiter_io_slave_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiArbiter_io_slave_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiArbiter_io_slave_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiArbiter_io_slave_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiArbiter_io_slave_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiArbiter_io_slave_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiArbiter_io_slave_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiArbiter_io_slave_aw_valid;
  assign io_slaves_1_r_ready = NastiArbiter_1_io_slave_r_ready;
  assign io_slaves_1_ar_bits_user = NastiArbiter_1_io_slave_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiArbiter_1_io_slave_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiArbiter_1_io_slave_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiArbiter_1_io_slave_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiArbiter_1_io_slave_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiArbiter_1_io_slave_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiArbiter_1_io_slave_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiArbiter_1_io_slave_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiArbiter_1_io_slave_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiArbiter_1_io_slave_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiArbiter_1_io_slave_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiArbiter_1_io_slave_ar_valid;
  assign io_slaves_1_b_ready = NastiArbiter_1_io_slave_b_ready;
  assign io_slaves_1_w_bits_user = NastiArbiter_1_io_slave_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiArbiter_1_io_slave_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiArbiter_1_io_slave_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiArbiter_1_io_slave_w_bits_data;
  assign io_slaves_1_w_valid = NastiArbiter_1_io_slave_w_valid;
  assign io_slaves_1_aw_bits_user = NastiArbiter_1_io_slave_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiArbiter_1_io_slave_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiArbiter_1_io_slave_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiArbiter_1_io_slave_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiArbiter_1_io_slave_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiArbiter_1_io_slave_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiArbiter_1_io_slave_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiArbiter_1_io_slave_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiArbiter_1_io_slave_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiArbiter_1_io_slave_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiArbiter_1_io_slave_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiArbiter_1_io_slave_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  assign io_masters_1_r_bits_user = NastiRouter_1_io_master_r_bits_user;
  assign io_masters_1_r_bits_id = NastiRouter_1_io_master_r_bits_id;
  assign io_masters_1_r_bits_last = NastiRouter_1_io_master_r_bits_last;
  assign io_masters_1_r_bits_data = NastiRouter_1_io_master_r_bits_data;
  assign io_masters_1_r_bits_resp = NastiRouter_1_io_master_r_bits_resp;
  assign io_masters_1_r_valid = NastiRouter_1_io_master_r_valid;
  assign io_masters_1_ar_ready = NastiRouter_1_io_master_ar_ready;
  assign io_masters_1_b_bits_user = NastiRouter_1_io_master_b_bits_user;
  assign io_masters_1_b_bits_id = NastiRouter_1_io_master_b_bits_id;
  assign io_masters_1_b_bits_resp = NastiRouter_1_io_master_b_bits_resp;
  assign io_masters_1_b_valid = NastiRouter_1_io_master_b_valid;
  assign io_masters_1_w_ready = NastiRouter_1_io_master_w_ready;
  assign io_masters_1_aw_ready = NastiRouter_1_io_master_aw_ready;
  NastiRouter_0 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user )
  );
  NastiRouter_0 NastiRouter_1(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_1_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_1_aw_valid ),
       .io_master_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_master_w_ready( NastiRouter_1_io_master_w_ready ),
       .io_master_w_valid( io_masters_1_w_valid ),
       .io_master_w_bits_data( io_masters_1_w_bits_data ),
       .io_master_w_bits_last( io_masters_1_w_bits_last ),
       .io_master_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_master_w_bits_user( io_masters_1_w_bits_user ),
       .io_master_b_ready( io_masters_1_b_ready ),
       .io_master_b_valid( NastiRouter_1_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_1_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_1_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_1_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_1_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_1_ar_valid ),
       .io_master_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_master_r_ready( io_masters_1_r_ready ),
       .io_master_r_valid( NastiRouter_1_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_1_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_1_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_1_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_1_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_1_io_master_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_slave_0_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_1_r_bits_user )
  );
  NastiArbiter_1 NastiArbiter(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_master_1_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_master_1_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_master_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_master_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_0_w_ready ),
       .io_slave_w_valid( NastiArbiter_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_0_b_valid ),
       .io_slave_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_0_r_valid ),
       .io_slave_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiArbiter_1 NastiArbiter_1(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_master_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_master_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_master_0_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_master_0_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_1_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_1_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_1_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_1_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_1_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_1_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_1_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_1_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_1_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_1_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_1_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_1_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_1_w_ready ),
       .io_slave_w_valid( NastiArbiter_1_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_1_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_1_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_1_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_1_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_1_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_1_b_valid ),
       .io_slave_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_1_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_1_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_1_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_1_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_1_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_1_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_1_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_1_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_1_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_1_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_1_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_1_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_1_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_1_r_valid ),
       .io_slave_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_1_r_bits_user )
  );
endmodule

module RRArbiter_6(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [5:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [5:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [5:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [5:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[5:0] io_out_bits_id,
    output io_out_bits_user,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg [1:0] last_grant;
  wire[1:0] T89;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire T22;
  wire[5:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T11 ? 2'h1 : T0;
  assign T0 = T9 ? 2'h2 : T1;
  assign T1 = T5 ? 2'h3 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : T4;
  assign T4 = io_in_2_valid ? 2'h2 : 2'h3;
  assign T5 = io_in_3_valid & T6;
  assign T6 = last_grant < 2'h3;
  assign T89 = reset ? 2'h0 : T7;
  assign T7 = T8 ? chosen : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_2_valid & T10;
  assign T10 = last_grant < 2'h2;
  assign T11 = io_in_1_valid & T12;
  assign T12 = last_grant < 2'h1;
  assign io_out_bits_user = T13;
  assign T13 = T19 ? T17 : T14;
  assign T14 = T15 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T15 = T16[1'h0];
  assign T16 = chosen;
  assign T17 = T18 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T18 = T16[1'h0];
  assign T19 = T16[1'h1];
  assign io_out_bits_id = T20;
  assign T20 = T25 ? T23 : T21;
  assign T21 = T22 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T22 = T16[1'h0];
  assign T23 = T24 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T24 = T16[1'h0];
  assign T25 = T16[1'h1];
  assign io_out_bits_resp = T26;
  assign T26 = T31 ? T29 : T27;
  assign T27 = T28 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T28 = T16[1'h0];
  assign T29 = T30 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T30 = T16[1'h0];
  assign T31 = T16[1'h1];
  assign io_out_valid = T32;
  assign T32 = T37 ? T35 : T33;
  assign T33 = T34 ? io_in_1_valid : io_in_0_valid;
  assign T34 = T16[1'h0];
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T16[1'h0];
  assign T37 = T16[1'h1];
  assign io_in_0_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T52 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T44 | T42;
  assign T42 = io_in_3_valid & T43;
  assign T43 = last_grant < 2'h3;
  assign T44 = T47 | T45;
  assign T45 = io_in_2_valid & T46;
  assign T46 = last_grant < 2'h2;
  assign T47 = T50 | T48;
  assign T48 = io_in_1_valid & T49;
  assign T49 = last_grant < 2'h1;
  assign T50 = io_in_0_valid & T51;
  assign T51 = last_grant < 2'h0;
  assign T52 = last_grant < 2'h0;
  assign io_in_1_ready = T53;
  assign T53 = T54 & io_out_ready;
  assign T54 = T60 | T55;
  assign T55 = T56 ^ 1'h1;
  assign T56 = T57 | io_in_0_valid;
  assign T57 = T58 | T42;
  assign T58 = T59 | T45;
  assign T59 = T50 | T48;
  assign T60 = T62 & T61;
  assign T61 = last_grant < 2'h1;
  assign T62 = T50 ^ 1'h1;
  assign io_in_2_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T71 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_1_valid;
  assign T67 = T68 | io_in_0_valid;
  assign T68 = T69 | T42;
  assign T69 = T70 | T45;
  assign T70 = T50 | T48;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T50 | T48;
  assign io_in_3_ready = T75;
  assign T75 = T76 & io_out_ready;
  assign T76 = T84 | T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T79 | io_in_2_valid;
  assign T79 = T80 | io_in_1_valid;
  assign T80 = T81 | io_in_0_valid;
  assign T81 = T82 | T42;
  assign T82 = T83 | T45;
  assign T83 = T50 | T48;
  assign T84 = T86 & T85;
  assign T85 = last_grant < 2'h3;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | T45;
  assign T88 = T50 | T48;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= chosen;
    end
  end
endmodule

module JunctionsPeekingArbiter_1(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [63:0] io_in_3_bits_data,
    input  io_in_3_bits_last,
    input [5:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [63:0] io_in_2_bits_data,
    input  io_in_2_bits_last,
    input [5:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_last,
    input [5:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_last,
    input [5:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[63:0] io_out_bits_data,
    output io_out_bits_last,
    output[5:0] io_out_bits_id,
    output io_out_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] chosen;
  wire[1:0] choice;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  reg [1:0] T7;
  wire[1:0] T9;
  wire[1:0] T10;
  reg [1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  reg [1:0] T15;
  wire[1:0] T16;
  reg [1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  reg [1:0] T40;
  wire[1:0] T41;
  reg [1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  reg [1:0] T64;
  wire[1:0] T135;
  wire[2:0] T65;
  wire[2:0] T136;
  reg [1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[2:0] T137;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T138;
  wire[2:0] T74;
  wire[2:0] T139;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[2:0] T140;
  reg [1:0] lockIdx;
  wire[1:0] T141;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire T90;
  reg  locked;
  wire T142;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[5:0] T97;
  wire[5:0] T98;
  wire T99;
  wire[5:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[63:0] T109;
  wire[63:0] T110;
  wire T111;
  wire[63:0] T112;
  wire T113;
  wire T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_user = T0;
  assign T0 = T96 ? T94 : T1;
  assign T1 = T2 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T2 = T3[1'h0];
  assign T3 = chosen;
  assign chosen = locked ? lockIdx : choice;
  assign choice = T69 ? T63 : T4;
  assign T4 = T45 ? T39 : T5;
  assign T5 = T20 ? T14 : T6;
  assign T6 = T13 ? T11 : T7;
  always @(*) case (T9)
    0: T7 = 2'h0;
    1: T7 = 2'h1;
    2: T7 = 2'h2;
    3: T7 = 2'h3;
    default: begin
      T7 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T7 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T9 = T10 - 2'h1;
  assign T10 = lockIdx + 2'h1;
  always @(*) case (T12)
    0: T11 = 2'h0;
    1: T11 = 2'h1;
    2: T11 = 2'h2;
    3: T11 = 2'h3;
    default: begin
      T11 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T11 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T12 = 2'h3 + T10;
  assign T13 = T10 < 2'h1;
  assign T14 = T19 ? T17 : T15;
  always @(*) case (T16)
    0: T15 = 2'h0;
    1: T15 = 2'h1;
    2: T15 = 2'h2;
    3: T15 = 2'h3;
    default: begin
      T15 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T15 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T16 = T10 - 2'h2;
  always @(*) case (T18)
    0: T17 = 2'h0;
    1: T17 = 2'h1;
    2: T17 = 2'h2;
    3: T17 = 2'h3;
    default: begin
      T17 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T17 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T18 = 2'h2 + T10;
  assign T19 = T10 < 2'h2;
  assign T20 = T38 ? T30 : T21;
  assign T21 = T29 ? T27 : T22;
  assign T22 = T23 ? io_in_1_valid : io_in_0_valid;
  assign T23 = T24[1'h0];
  assign T24 = T25;
  assign T25 = T26 - 2'h2;
  assign T26 = lockIdx + 2'h1;
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T24[1'h0];
  assign T29 = T24[1'h1];
  assign T30 = T37 ? T35 : T31;
  assign T31 = T32 ? io_in_1_valid : io_in_0_valid;
  assign T32 = T33[1'h0];
  assign T33 = T34;
  assign T34 = 2'h2 + T26;
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T33[1'h0];
  assign T37 = T33[1'h1];
  assign T38 = T26 < 2'h2;
  assign T39 = T44 ? T42 : T40;
  always @(*) case (T41)
    0: T40 = 2'h0;
    1: T40 = 2'h1;
    2: T40 = 2'h2;
    3: T40 = 2'h3;
    default: begin
      T40 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T40 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T41 = T10 - 2'h3;
  always @(*) case (T43)
    0: T42 = 2'h0;
    1: T42 = 2'h1;
    2: T42 = 2'h2;
    3: T42 = 2'h3;
    default: begin
      T42 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T42 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T43 = 2'h1 + T10;
  assign T44 = T10 < 2'h3;
  assign T45 = T62 ? T54 : T46;
  assign T46 = T53 ? T51 : T47;
  assign T47 = T48 ? io_in_1_valid : io_in_0_valid;
  assign T48 = T49[1'h0];
  assign T49 = T50;
  assign T50 = T26 - 2'h3;
  assign T51 = T52 ? io_in_3_valid : io_in_2_valid;
  assign T52 = T49[1'h0];
  assign T53 = T49[1'h1];
  assign T54 = T61 ? T59 : T55;
  assign T55 = T56 ? io_in_1_valid : io_in_0_valid;
  assign T56 = T57[1'h0];
  assign T57 = T58;
  assign T58 = 2'h1 + T26;
  assign T59 = T60 ? io_in_3_valid : io_in_2_valid;
  assign T60 = T57[1'h0];
  assign T61 = T57[1'h1];
  assign T62 = T26 < 2'h3;
  assign T63 = T68 ? T66 : T64;
  always @(*) case (T135)
    0: T64 = 2'h0;
    1: T64 = 2'h1;
    2: T64 = 2'h2;
    3: T64 = 2'h3;
    default: begin
      T64 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T64 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T135 = T65[1'h1:1'h0];
  assign T65 = T136 - 3'h4;
  assign T136 = {1'h0, T10};
  always @(*) case (T67)
    0: T66 = 2'h0;
    1: T66 = 2'h1;
    2: T66 = 2'h2;
    3: T66 = 2'h3;
    default: begin
      T66 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T66 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T67 = 2'h0 + T10;
  assign T68 = T137 < 3'h4;
  assign T137 = {1'h0, T10};
  assign T69 = T86 ? T78 : T70;
  assign T70 = T77 ? T75 : T71;
  assign T71 = T72 ? io_in_1_valid : io_in_0_valid;
  assign T72 = T73[1'h0];
  assign T73 = T138;
  assign T138 = T74[1'h1:1'h0];
  assign T74 = T139 - 3'h4;
  assign T139 = {1'h0, T26};
  assign T75 = T76 ? io_in_3_valid : io_in_2_valid;
  assign T76 = T73[1'h0];
  assign T77 = T73[1'h1];
  assign T78 = T85 ? T83 : T79;
  assign T79 = T80 ? io_in_1_valid : io_in_0_valid;
  assign T80 = T81[1'h0];
  assign T81 = T82;
  assign T82 = 2'h0 + T26;
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T81[1'h0];
  assign T85 = T81[1'h1];
  assign T86 = T140 < 3'h4;
  assign T140 = {1'h0, T26};
  assign T141 = reset ? 2'h0 : T87;
  assign T87 = T88 ? choice : lockIdx;
  assign T88 = T90 & T89;
  assign T89 = locked ^ 1'h1;
  assign T90 = io_out_ready & io_out_valid;
  assign T142 = reset ? 1'h0 : T91;
  assign T91 = T93 ? 1'h0 : T92;
  assign T92 = T88 ? 1'h1 : locked;
  assign T93 = T90 & io_out_bits_last;
  assign T94 = T95 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T95 = T3[1'h0];
  assign T96 = T3[1'h1];
  assign io_out_bits_id = T97;
  assign T97 = T102 ? T100 : T98;
  assign T98 = T99 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T99 = T3[1'h0];
  assign T100 = T101 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T101 = T3[1'h0];
  assign T102 = T3[1'h1];
  assign io_out_bits_last = T103;
  assign T103 = T108 ? T106 : T104;
  assign T104 = T105 ? io_in_1_bits_last : io_in_0_bits_last;
  assign T105 = T3[1'h0];
  assign T106 = T107 ? io_in_3_bits_last : io_in_2_bits_last;
  assign T107 = T3[1'h0];
  assign T108 = T3[1'h1];
  assign io_out_bits_data = T109;
  assign T109 = T114 ? T112 : T110;
  assign T110 = T111 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T111 = T3[1'h0];
  assign T112 = T113 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T113 = T3[1'h0];
  assign T114 = T3[1'h1];
  assign io_out_bits_resp = T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T117 = T3[1'h0];
  assign T118 = T119 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T119 = T3[1'h0];
  assign T120 = T3[1'h1];
  assign io_out_valid = T121;
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? io_in_1_valid : io_in_0_valid;
  assign T123 = T3[1'h0];
  assign T124 = T125 ? io_in_3_valid : io_in_2_valid;
  assign T125 = T3[1'h0];
  assign T126 = T3[1'h1];
  assign io_in_0_ready = T127;
  assign T127 = io_out_ready & T128;
  assign T128 = chosen == 2'h0;
  assign io_in_1_ready = T129;
  assign T129 = io_out_ready & T130;
  assign T130 = chosen == 2'h1;
  assign io_in_2_ready = T131;
  assign T131 = io_out_ready & T132;
  assign T132 = chosen == 2'h2;
  assign io_in_3_ready = T133;
  assign T133 = io_out_ready & T134;
  assign T134 = chosen == 2'h3;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h0;
    end else if(T88) begin
      lockIdx <= choice;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T93) begin
      locked <= 1'h0;
    end else if(T88) begin
      locked <= 1'h1;
    end
  end
endmodule

module NastiRouter_1(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [5:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[5:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [5:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[5:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_2_aw_ready,
    output io_slave_2_aw_valid,
    output[31:0] io_slave_2_aw_bits_addr,
    output[7:0] io_slave_2_aw_bits_len,
    output[2:0] io_slave_2_aw_bits_size,
    output[1:0] io_slave_2_aw_bits_burst,
    output io_slave_2_aw_bits_lock,
    output[3:0] io_slave_2_aw_bits_cache,
    output[2:0] io_slave_2_aw_bits_prot,
    output[3:0] io_slave_2_aw_bits_qos,
    output[3:0] io_slave_2_aw_bits_region,
    output[5:0] io_slave_2_aw_bits_id,
    output io_slave_2_aw_bits_user,
    input  io_slave_2_w_ready,
    output io_slave_2_w_valid,
    output[63:0] io_slave_2_w_bits_data,
    output io_slave_2_w_bits_last,
    output[7:0] io_slave_2_w_bits_strb,
    output io_slave_2_w_bits_user,
    output io_slave_2_b_ready,
    input  io_slave_2_b_valid,
    input [1:0] io_slave_2_b_bits_resp,
    input [5:0] io_slave_2_b_bits_id,
    input  io_slave_2_b_bits_user,
    input  io_slave_2_ar_ready,
    output io_slave_2_ar_valid,
    output[31:0] io_slave_2_ar_bits_addr,
    output[7:0] io_slave_2_ar_bits_len,
    output[2:0] io_slave_2_ar_bits_size,
    output[1:0] io_slave_2_ar_bits_burst,
    output io_slave_2_ar_bits_lock,
    output[3:0] io_slave_2_ar_bits_cache,
    output[2:0] io_slave_2_ar_bits_prot,
    output[3:0] io_slave_2_ar_bits_qos,
    output[3:0] io_slave_2_ar_bits_region,
    output[5:0] io_slave_2_ar_bits_id,
    output io_slave_2_ar_bits_user,
    output io_slave_2_r_ready,
    input  io_slave_2_r_valid,
    input [1:0] io_slave_2_r_bits_resp,
    input [63:0] io_slave_2_r_bits_data,
    input  io_slave_2_r_bits_last,
    input [5:0] io_slave_2_r_bits_id,
    input  io_slave_2_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[5:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [5:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[5:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [5:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[5:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [5:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[5:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [5:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[2:0] ar_route;
  wire[2:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire w_invalid;
  wire T14;
  wire[2:0] aw_route;
  wire[2:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T82;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg  R40;
  wire T83;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  R51;
  wire T84;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire ar_ready;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire w_ready;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire aw_ready;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire b_arb_io_in_3_ready;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[5:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_3_ready;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[5:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[5:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[5:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R29 = {1{$random}};
    R40 = {1{$random}};
    R51 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 3'h0;
  assign ar_route = T2;
  assign T2 = {T10, T3};
  assign T3 = {T7, T4};
  assign T4 = T6 & T5;
  assign T5 = io_master_ar_bits_addr < 32'h40008000;
  assign T6 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T7 = T9 & T8;
  assign T8 = io_master_ar_bits_addr < 32'h40010000;
  assign T9 = 32'h40008000 <= io_master_ar_bits_addr;
  assign T10 = T12 & T11;
  assign T11 = io_master_ar_bits_addr < 32'h40010200;
  assign T12 = 32'h40010000 <= io_master_ar_bits_addr;
  assign T13 = w_invalid & io_master_aw_valid;
  assign w_invalid = T14 ^ 1'h1;
  assign T14 = aw_route != 3'h0;
  assign aw_route = T15;
  assign T15 = {T23, T16};
  assign T16 = {T20, T17};
  assign T17 = T19 & T18;
  assign T18 = io_master_aw_bits_addr < 32'h40008000;
  assign T19 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T20 = T22 & T21;
  assign T21 = io_master_aw_bits_addr < 32'h40010000;
  assign T22 = 32'h40008000 <= io_master_aw_bits_addr;
  assign T23 = T25 & T24;
  assign T24 = io_master_aw_bits_addr < 32'h40010200;
  assign T25 = 32'h40010000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T26;
  assign T26 = io_master_ar_valid & T27;
  assign T27 = ar_route[1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T28;
  assign T28 = io_master_w_valid & R29;
  assign T82 = reset ? 1'h0 : T30;
  assign T30 = T33 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : R29;
  assign T32 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T33 = T34 & io_slave_0_w_bits_last;
  assign T34 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T35;
  assign T35 = io_master_aw_valid & T36;
  assign T36 = aw_route[1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T37;
  assign T37 = io_master_ar_valid & T38;
  assign T38 = ar_route[1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T39;
  assign T39 = io_master_w_valid & R40;
  assign T83 = reset ? 1'h0 : T41;
  assign T41 = T44 ? 1'h0 : T42;
  assign T42 = T43 ? 1'h1 : R40;
  assign T43 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T44 = T45 & io_slave_1_w_bits_last;
  assign T45 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T46;
  assign T46 = io_master_aw_valid & T47;
  assign T47 = aw_route[1'h1];
  assign io_slave_2_r_ready = r_arb_io_in_2_ready;
  assign io_slave_2_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_2_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_2_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_2_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_2_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_2_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_2_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_2_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_2_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_2_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_2_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_2_ar_valid = T48;
  assign T48 = io_master_ar_valid & T49;
  assign T49 = ar_route[2'h2];
  assign io_slave_2_b_ready = b_arb_io_in_2_ready;
  assign io_slave_2_w_bits_user = io_master_w_bits_user;
  assign io_slave_2_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_2_w_bits_last = io_master_w_bits_last;
  assign io_slave_2_w_bits_data = io_master_w_bits_data;
  assign io_slave_2_w_valid = T50;
  assign T50 = io_master_w_valid & R51;
  assign T84 = reset ? 1'h0 : T52;
  assign T52 = T55 ? 1'h0 : T53;
  assign T53 = T54 ? 1'h1 : R51;
  assign T54 = io_slave_2_aw_ready & io_slave_2_aw_valid;
  assign T55 = T56 & io_slave_2_w_bits_last;
  assign T56 = io_slave_2_w_ready & io_slave_2_w_valid;
  assign io_slave_2_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_2_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_2_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_2_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_2_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_2_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_2_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_2_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_2_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_2_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_2_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_2_aw_valid = T57;
  assign T57 = io_master_aw_valid & T58;
  assign T58 = aw_route[2'h2];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T59;
  assign T59 = ar_ready | T60;
  assign T60 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T63 | T61;
  assign T61 = io_slave_2_ar_ready & T62;
  assign T62 = ar_route[2'h2];
  assign T63 = T66 | T64;
  assign T64 = io_slave_1_ar_ready & T65;
  assign T65 = ar_route[1'h1];
  assign T66 = io_slave_0_ar_ready & T67;
  assign T67 = ar_route[1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T68;
  assign T68 = w_ready | err_slave_io_w_ready;
  assign w_ready = T70 | T69;
  assign T69 = io_slave_2_w_ready & R51;
  assign T70 = T72 | T71;
  assign T71 = io_slave_1_w_ready & R40;
  assign T72 = io_slave_0_w_ready & R29;
  assign io_master_aw_ready = T73;
  assign T73 = aw_ready | T74;
  assign T74 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T77 | T75;
  assign T75 = io_slave_2_aw_ready & T76;
  assign T76 = aw_route[2'h2];
  assign T77 = T80 | T78;
  assign T78 = io_slave_1_aw_ready & T79;
  assign T79 = aw_route[1'h1];
  assign T80 = io_slave_0_aw_ready & T81;
  assign T81 = aw_route[1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T13 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_3_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_3_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_6 b_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( b_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_b_valid ),
       .io_in_3_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_3_bits_id( err_slave_io_b_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_b_valid ),
       .io_in_2_bits_resp( io_slave_2_b_bits_resp ),
       .io_in_2_bits_id( io_slave_2_b_bits_id ),
       .io_in_2_bits_user( io_slave_2_b_bits_user ),
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter_1 r_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( r_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_r_valid ),
       .io_in_3_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_3_bits_data( err_slave_io_r_bits_data ),
       .io_in_3_bits_last( err_slave_io_r_bits_last ),
       .io_in_3_bits_id( err_slave_io_r_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_r_valid ),
       .io_in_2_bits_resp( io_slave_2_r_bits_resp ),
       .io_in_2_bits_data( io_slave_2_r_bits_data ),
       .io_in_2_bits_last( io_slave_2_r_bits_last ),
       .io_in_2_bits_id( io_slave_2_r_bits_id ),
       .io_in_2_bits_user( io_slave_2_r_bits_user ),
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R29 <= 1'h0;
    end else if(T33) begin
      R29 <= 1'h0;
    end else if(T32) begin
      R29 <= 1'h1;
    end
    if(reset) begin
      R40 <= 1'h0;
    end else if(T44) begin
      R40 <= 1'h0;
    end else if(T43) begin
      R40 <= 1'h1;
    end
    if(reset) begin
      R51 <= 1'h0;
    end else if(T55) begin
      R51 <= 1'h0;
    end else if(T54) begin
      R51 <= 1'h1;
    end
  end
endmodule

module NastiCrossbar_1(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [5:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[5:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [5:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[5:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[5:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [5:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[5:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [5:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[5:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [5:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[5:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [5:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[5:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [5:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[5:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [5:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[5:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[5:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_2_aw_bits_burst;
  wire NastiRouter_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_region;
  wire[5:0] NastiRouter_io_slave_2_aw_bits_id;
  wire NastiRouter_io_slave_2_aw_bits_user;
  wire NastiRouter_io_slave_2_w_valid;
  wire[63:0] NastiRouter_io_slave_2_w_bits_data;
  wire NastiRouter_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_io_slave_2_w_bits_strb;
  wire NastiRouter_io_slave_2_w_bits_user;
  wire NastiRouter_io_slave_2_b_ready;
  wire NastiRouter_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_2_ar_bits_burst;
  wire NastiRouter_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_region;
  wire[5:0] NastiRouter_io_slave_2_ar_bits_id;
  wire NastiRouter_io_slave_2_ar_bits_user;
  wire NastiRouter_io_slave_2_r_ready;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[5:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[5:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[5:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[5:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiRouter_io_slave_0_r_ready;
  assign io_slaves_0_ar_bits_user = NastiRouter_io_slave_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiRouter_io_slave_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiRouter_io_slave_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiRouter_io_slave_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiRouter_io_slave_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiRouter_io_slave_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiRouter_io_slave_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiRouter_io_slave_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiRouter_io_slave_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiRouter_io_slave_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiRouter_io_slave_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiRouter_io_slave_0_ar_valid;
  assign io_slaves_0_b_ready = NastiRouter_io_slave_0_b_ready;
  assign io_slaves_0_w_bits_user = NastiRouter_io_slave_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiRouter_io_slave_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiRouter_io_slave_0_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiRouter_io_slave_0_w_bits_data;
  assign io_slaves_0_w_valid = NastiRouter_io_slave_0_w_valid;
  assign io_slaves_0_aw_bits_user = NastiRouter_io_slave_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiRouter_io_slave_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiRouter_io_slave_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiRouter_io_slave_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiRouter_io_slave_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiRouter_io_slave_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiRouter_io_slave_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiRouter_io_slave_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiRouter_io_slave_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiRouter_io_slave_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiRouter_io_slave_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiRouter_io_slave_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRouter_io_slave_1_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRouter_io_slave_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRouter_io_slave_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRouter_io_slave_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRouter_io_slave_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRouter_io_slave_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRouter_io_slave_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRouter_io_slave_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRouter_io_slave_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRouter_io_slave_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRouter_io_slave_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRouter_io_slave_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRouter_io_slave_1_ar_valid;
  assign io_slaves_1_b_ready = NastiRouter_io_slave_1_b_ready;
  assign io_slaves_1_w_bits_user = NastiRouter_io_slave_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRouter_io_slave_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRouter_io_slave_1_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRouter_io_slave_1_w_bits_data;
  assign io_slaves_1_w_valid = NastiRouter_io_slave_1_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRouter_io_slave_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRouter_io_slave_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRouter_io_slave_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRouter_io_slave_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRouter_io_slave_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRouter_io_slave_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRouter_io_slave_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRouter_io_slave_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRouter_io_slave_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRouter_io_slave_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRouter_io_slave_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRouter_io_slave_1_aw_valid;
  assign io_slaves_2_r_ready = NastiRouter_io_slave_2_r_ready;
  assign io_slaves_2_ar_bits_user = NastiRouter_io_slave_2_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiRouter_io_slave_2_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiRouter_io_slave_2_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiRouter_io_slave_2_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiRouter_io_slave_2_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiRouter_io_slave_2_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiRouter_io_slave_2_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiRouter_io_slave_2_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiRouter_io_slave_2_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiRouter_io_slave_2_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiRouter_io_slave_2_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiRouter_io_slave_2_ar_valid;
  assign io_slaves_2_b_ready = NastiRouter_io_slave_2_b_ready;
  assign io_slaves_2_w_bits_user = NastiRouter_io_slave_2_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiRouter_io_slave_2_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiRouter_io_slave_2_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiRouter_io_slave_2_w_bits_data;
  assign io_slaves_2_w_valid = NastiRouter_io_slave_2_w_valid;
  assign io_slaves_2_aw_bits_user = NastiRouter_io_slave_2_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiRouter_io_slave_2_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiRouter_io_slave_2_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiRouter_io_slave_2_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiRouter_io_slave_2_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiRouter_io_slave_2_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiRouter_io_slave_2_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiRouter_io_slave_2_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiRouter_io_slave_2_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiRouter_io_slave_2_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiRouter_io_slave_2_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiRouter_io_slave_2_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  NastiRouter_1 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_2_aw_ready( io_slaves_2_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( io_slaves_2_w_ready ),
       .io_slave_2_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_slave_2_b_valid( io_slaves_2_b_valid ),
       .io_slave_2_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slave_2_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slave_2_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slave_2_ar_ready( io_slaves_2_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_slave_2_r_valid( io_slaves_2_r_valid ),
       .io_slave_2_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slave_2_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slave_2_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slave_2_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slave_2_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slave_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( io_slaves_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( io_slaves_1_b_valid ),
       .io_slave_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( io_slaves_1_r_valid ),
       .io_slave_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slave_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( io_slaves_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( io_slaves_0_b_valid ),
       .io_slave_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( io_slaves_0_r_valid ),
       .io_slave_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [5:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[5:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [5:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[5:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[5:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [5:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[5:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [5:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[5:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [5:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[5:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [5:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[5:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [5:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[5:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [5:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[5:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[5:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_2_aw_valid;
  wire[31:0] xbar_io_slaves_2_aw_bits_addr;
  wire[7:0] xbar_io_slaves_2_aw_bits_len;
  wire[2:0] xbar_io_slaves_2_aw_bits_size;
  wire[1:0] xbar_io_slaves_2_aw_bits_burst;
  wire xbar_io_slaves_2_aw_bits_lock;
  wire[3:0] xbar_io_slaves_2_aw_bits_cache;
  wire[2:0] xbar_io_slaves_2_aw_bits_prot;
  wire[3:0] xbar_io_slaves_2_aw_bits_qos;
  wire[3:0] xbar_io_slaves_2_aw_bits_region;
  wire[5:0] xbar_io_slaves_2_aw_bits_id;
  wire xbar_io_slaves_2_aw_bits_user;
  wire xbar_io_slaves_2_w_valid;
  wire[63:0] xbar_io_slaves_2_w_bits_data;
  wire xbar_io_slaves_2_w_bits_last;
  wire[7:0] xbar_io_slaves_2_w_bits_strb;
  wire xbar_io_slaves_2_w_bits_user;
  wire xbar_io_slaves_2_b_ready;
  wire xbar_io_slaves_2_ar_valid;
  wire[31:0] xbar_io_slaves_2_ar_bits_addr;
  wire[7:0] xbar_io_slaves_2_ar_bits_len;
  wire[2:0] xbar_io_slaves_2_ar_bits_size;
  wire[1:0] xbar_io_slaves_2_ar_bits_burst;
  wire xbar_io_slaves_2_ar_bits_lock;
  wire[3:0] xbar_io_slaves_2_ar_bits_cache;
  wire[2:0] xbar_io_slaves_2_ar_bits_prot;
  wire[3:0] xbar_io_slaves_2_ar_bits_qos;
  wire[3:0] xbar_io_slaves_2_ar_bits_region;
  wire[5:0] xbar_io_slaves_2_ar_bits_id;
  wire xbar_io_slaves_2_ar_bits_user;
  wire xbar_io_slaves_2_r_ready;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[5:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[5:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[5:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[5:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = xbar_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = xbar_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = xbar_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = xbar_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = xbar_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = xbar_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = xbar_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = xbar_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = xbar_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = xbar_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = xbar_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = xbar_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = xbar_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = xbar_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = xbar_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = xbar_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = xbar_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = xbar_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = xbar_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = xbar_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = xbar_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = xbar_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = xbar_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = xbar_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = xbar_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = xbar_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = xbar_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = xbar_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = xbar_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = xbar_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = xbar_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = xbar_io_slaves_1_r_ready;
  assign io_slaves_1_ar_bits_user = xbar_io_slaves_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = xbar_io_slaves_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = xbar_io_slaves_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = xbar_io_slaves_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = xbar_io_slaves_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = xbar_io_slaves_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = xbar_io_slaves_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = xbar_io_slaves_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = xbar_io_slaves_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = xbar_io_slaves_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = xbar_io_slaves_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = xbar_io_slaves_1_ar_valid;
  assign io_slaves_1_b_ready = xbar_io_slaves_1_b_ready;
  assign io_slaves_1_w_bits_user = xbar_io_slaves_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = xbar_io_slaves_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = xbar_io_slaves_1_w_bits_last;
  assign io_slaves_1_w_bits_data = xbar_io_slaves_1_w_bits_data;
  assign io_slaves_1_w_valid = xbar_io_slaves_1_w_valid;
  assign io_slaves_1_aw_bits_user = xbar_io_slaves_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = xbar_io_slaves_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = xbar_io_slaves_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = xbar_io_slaves_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = xbar_io_slaves_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = xbar_io_slaves_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = xbar_io_slaves_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = xbar_io_slaves_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = xbar_io_slaves_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = xbar_io_slaves_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = xbar_io_slaves_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = xbar_io_slaves_1_aw_valid;
  assign io_slaves_2_r_ready = xbar_io_slaves_2_r_ready;
  assign io_slaves_2_ar_bits_user = xbar_io_slaves_2_ar_bits_user;
  assign io_slaves_2_ar_bits_id = xbar_io_slaves_2_ar_bits_id;
  assign io_slaves_2_ar_bits_region = xbar_io_slaves_2_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = xbar_io_slaves_2_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = xbar_io_slaves_2_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = xbar_io_slaves_2_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = xbar_io_slaves_2_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = xbar_io_slaves_2_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = xbar_io_slaves_2_ar_bits_size;
  assign io_slaves_2_ar_bits_len = xbar_io_slaves_2_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = xbar_io_slaves_2_ar_bits_addr;
  assign io_slaves_2_ar_valid = xbar_io_slaves_2_ar_valid;
  assign io_slaves_2_b_ready = xbar_io_slaves_2_b_ready;
  assign io_slaves_2_w_bits_user = xbar_io_slaves_2_w_bits_user;
  assign io_slaves_2_w_bits_strb = xbar_io_slaves_2_w_bits_strb;
  assign io_slaves_2_w_bits_last = xbar_io_slaves_2_w_bits_last;
  assign io_slaves_2_w_bits_data = xbar_io_slaves_2_w_bits_data;
  assign io_slaves_2_w_valid = xbar_io_slaves_2_w_valid;
  assign io_slaves_2_aw_bits_user = xbar_io_slaves_2_aw_bits_user;
  assign io_slaves_2_aw_bits_id = xbar_io_slaves_2_aw_bits_id;
  assign io_slaves_2_aw_bits_region = xbar_io_slaves_2_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = xbar_io_slaves_2_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = xbar_io_slaves_2_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = xbar_io_slaves_2_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = xbar_io_slaves_2_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = xbar_io_slaves_2_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = xbar_io_slaves_2_aw_bits_size;
  assign io_slaves_2_aw_bits_len = xbar_io_slaves_2_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = xbar_io_slaves_2_aw_bits_addr;
  assign io_slaves_2_aw_valid = xbar_io_slaves_2_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  NastiCrossbar_1 xbar(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_2_aw_ready ),
       .io_slaves_2_aw_valid( xbar_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( xbar_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( xbar_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( xbar_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( xbar_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( xbar_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( xbar_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( xbar_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( xbar_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( xbar_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( xbar_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( xbar_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_2_w_ready ),
       .io_slaves_2_w_valid( xbar_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( xbar_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( xbar_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( xbar_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( xbar_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( xbar_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_2_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_2_ar_ready ),
       .io_slaves_2_ar_valid( xbar_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( xbar_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( xbar_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( xbar_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( xbar_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( xbar_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( xbar_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( xbar_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( xbar_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( xbar_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( xbar_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( xbar_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( xbar_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_2_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_1_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_1_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_1_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect_1(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [5:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[5:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [5:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[5:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [5:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[5:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [5:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[5:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[5:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [5:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[5:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [5:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[5:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [5:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[5:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [5:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[5:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [5:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[5:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [5:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiErrorSlave_io_aw_ready;
  wire NastiErrorSlave_io_w_ready;
  wire NastiErrorSlave_io_b_valid;
  wire[1:0] NastiErrorSlave_io_b_bits_resp;
  wire[5:0] NastiErrorSlave_io_b_bits_id;
  wire NastiErrorSlave_io_ar_ready;
  wire NastiErrorSlave_io_r_valid;
  wire[1:0] NastiErrorSlave_io_r_bits_resp;
  wire[63:0] NastiErrorSlave_io_r_bits_data;
  wire NastiErrorSlave_io_r_bits_last;
  wire[5:0] NastiErrorSlave_io_r_bits_id;
  wire xbar_io_masters_1_aw_ready;
  wire xbar_io_masters_1_w_ready;
  wire xbar_io_masters_1_b_valid;
  wire[1:0] xbar_io_masters_1_b_bits_resp;
  wire[5:0] xbar_io_masters_1_b_bits_id;
  wire xbar_io_masters_1_b_bits_user;
  wire xbar_io_masters_1_ar_ready;
  wire xbar_io_masters_1_r_valid;
  wire[1:0] xbar_io_masters_1_r_bits_resp;
  wire[63:0] xbar_io_masters_1_r_bits_data;
  wire xbar_io_masters_1_r_bits_last;
  wire[5:0] xbar_io_masters_1_r_bits_id;
  wire xbar_io_masters_1_r_bits_user;
  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[5:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[5:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[5:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[5:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[5:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[5:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;
  wire NastiRecursiveInterconnect_io_masters_0_aw_ready;
  wire NastiRecursiveInterconnect_io_masters_0_w_ready;
  wire NastiRecursiveInterconnect_io_masters_0_b_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_b_bits_resp;
  wire[5:0] NastiRecursiveInterconnect_io_masters_0_b_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_b_bits_user;
  wire NastiRecursiveInterconnect_io_masters_0_ar_ready;
  wire NastiRecursiveInterconnect_io_masters_0_r_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_r_bits_resp;
  wire[63:0] NastiRecursiveInterconnect_io_masters_0_r_bits_data;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_last;
  wire[5:0] NastiRecursiveInterconnect_io_masters_0_r_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_2_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_2_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_2_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_r_ready;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_r_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  wire[5:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = NastiRecursiveInterconnect_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = NastiRecursiveInterconnect_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = NastiRecursiveInterconnect_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRecursiveInterconnect_io_slaves_1_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  assign io_slaves_1_b_ready = NastiRecursiveInterconnect_io_slaves_1_b_ready;
  assign io_slaves_1_w_bits_user = NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  assign io_slaves_1_w_valid = NastiRecursiveInterconnect_io_slaves_1_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  assign io_slaves_2_r_ready = NastiRecursiveInterconnect_io_slaves_2_r_ready;
  assign io_slaves_2_ar_bits_user = NastiRecursiveInterconnect_io_slaves_2_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiRecursiveInterconnect_io_slaves_2_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiRecursiveInterconnect_io_slaves_2_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiRecursiveInterconnect_io_slaves_2_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiRecursiveInterconnect_io_slaves_2_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiRecursiveInterconnect_io_slaves_2_ar_valid;
  assign io_slaves_2_b_ready = NastiRecursiveInterconnect_io_slaves_2_b_ready;
  assign io_slaves_2_w_bits_user = NastiRecursiveInterconnect_io_slaves_2_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiRecursiveInterconnect_io_slaves_2_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiRecursiveInterconnect_io_slaves_2_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiRecursiveInterconnect_io_slaves_2_w_bits_data;
  assign io_slaves_2_w_valid = NastiRecursiveInterconnect_io_slaves_2_w_valid;
  assign io_slaves_2_aw_bits_user = NastiRecursiveInterconnect_io_slaves_2_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiRecursiveInterconnect_io_slaves_2_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiRecursiveInterconnect_io_slaves_2_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiRecursiveInterconnect_io_slaves_2_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiRecursiveInterconnect_io_slaves_2_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiRecursiveInterconnect_io_slaves_2_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  assign io_masters_1_r_bits_user = xbar_io_masters_1_r_bits_user;
  assign io_masters_1_r_bits_id = xbar_io_masters_1_r_bits_id;
  assign io_masters_1_r_bits_last = xbar_io_masters_1_r_bits_last;
  assign io_masters_1_r_bits_data = xbar_io_masters_1_r_bits_data;
  assign io_masters_1_r_bits_resp = xbar_io_masters_1_r_bits_resp;
  assign io_masters_1_r_valid = xbar_io_masters_1_r_valid;
  assign io_masters_1_ar_ready = xbar_io_masters_1_ar_ready;
  assign io_masters_1_b_bits_user = xbar_io_masters_1_b_bits_user;
  assign io_masters_1_b_bits_id = xbar_io_masters_1_b_bits_id;
  assign io_masters_1_b_bits_resp = xbar_io_masters_1_b_bits_resp;
  assign io_masters_1_b_valid = xbar_io_masters_1_b_valid;
  assign io_masters_1_w_ready = xbar_io_masters_1_w_ready;
  assign io_masters_1_aw_ready = xbar_io_masters_1_aw_ready;
  NastiCrossbar_0 xbar(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( xbar_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( io_masters_1_aw_valid ),
       .io_masters_1_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_masters_1_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_masters_1_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_masters_1_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_masters_1_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_masters_1_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_masters_1_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_masters_1_w_ready( xbar_io_masters_1_w_ready ),
       .io_masters_1_w_valid( io_masters_1_w_valid ),
       .io_masters_1_w_bits_data( io_masters_1_w_bits_data ),
       .io_masters_1_w_bits_last( io_masters_1_w_bits_last ),
       .io_masters_1_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_masters_1_w_bits_user( io_masters_1_w_bits_user ),
       .io_masters_1_b_ready( io_masters_1_b_ready ),
       .io_masters_1_b_valid( xbar_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( xbar_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( xbar_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( xbar_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( xbar_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( io_masters_1_ar_valid ),
       .io_masters_1_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_masters_1_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_masters_1_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_masters_1_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_masters_1_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_masters_1_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_masters_1_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_masters_1_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_masters_1_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_masters_1_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_masters_1_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_masters_1_r_ready( io_masters_1_r_ready ),
       .io_masters_1_r_valid( xbar_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( xbar_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( xbar_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( xbar_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( xbar_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( xbar_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_1_aw_ready( NastiErrorSlave_io_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( NastiErrorSlave_io_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( NastiErrorSlave_io_b_valid ),
       .io_slaves_1_b_bits_resp( NastiErrorSlave_io_b_bits_resp ),
       .io_slaves_1_b_bits_id( NastiErrorSlave_io_b_bits_id ),
       //.io_slaves_1_b_bits_user(  )
       .io_slaves_1_ar_ready( NastiErrorSlave_io_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( NastiErrorSlave_io_r_valid ),
       .io_slaves_1_r_bits_resp( NastiErrorSlave_io_r_bits_resp ),
       .io_slaves_1_r_bits_data( NastiErrorSlave_io_r_bits_data ),
       .io_slaves_1_r_bits_last( NastiErrorSlave_io_r_bits_last ),
       .io_slaves_1_r_bits_id( NastiErrorSlave_io_r_bits_id ),
       //.io_slaves_1_r_bits_user(  )
       .io_slaves_0_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_slaves_0_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_slaves_0_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_slaves_0_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_slaves_0_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_slaves_0_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_slaves_0_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_slaves_0_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign xbar.io_slaves_1_b_bits_user = {1{$random}};
    assign xbar.io_slaves_1_r_bits_user = {1{$random}};
// synthesis translate_on
`endif
  NastiRecursiveInterconnect NastiRecursiveInterconnect(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_masters_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_masters_0_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_masters_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_masters_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_masters_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_masters_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_masters_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_masters_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_masters_0_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_masters_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_masters_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_masters_0_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_2_aw_ready ),
       .io_slaves_2_aw_valid( NastiRecursiveInterconnect_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( NastiRecursiveInterconnect_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( NastiRecursiveInterconnect_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( NastiRecursiveInterconnect_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( NastiRecursiveInterconnect_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( NastiRecursiveInterconnect_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_2_w_ready ),
       .io_slaves_2_w_valid( NastiRecursiveInterconnect_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( NastiRecursiveInterconnect_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( NastiRecursiveInterconnect_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( NastiRecursiveInterconnect_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( NastiRecursiveInterconnect_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( NastiRecursiveInterconnect_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_2_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_2_ar_ready ),
       .io_slaves_2_ar_valid( NastiRecursiveInterconnect_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( NastiRecursiveInterconnect_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( NastiRecursiveInterconnect_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( NastiRecursiveInterconnect_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( NastiRecursiveInterconnect_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( NastiRecursiveInterconnect_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( NastiRecursiveInterconnect_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_2_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_1_aw_valid( NastiRecursiveInterconnect_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( NastiRecursiveInterconnect_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( NastiRecursiveInterconnect_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( NastiRecursiveInterconnect_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( NastiRecursiveInterconnect_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( NastiRecursiveInterconnect_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_1_w_ready ),
       .io_slaves_1_w_valid( NastiRecursiveInterconnect_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( NastiRecursiveInterconnect_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( NastiRecursiveInterconnect_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( NastiRecursiveInterconnect_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( NastiRecursiveInterconnect_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( NastiRecursiveInterconnect_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_1_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_1_ar_valid( NastiRecursiveInterconnect_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( NastiRecursiveInterconnect_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( NastiRecursiveInterconnect_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( NastiRecursiveInterconnect_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( NastiRecursiveInterconnect_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( NastiRecursiveInterconnect_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( NastiRecursiveInterconnect_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_1_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( NastiRecursiveInterconnect_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( NastiRecursiveInterconnect_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( NastiRecursiveInterconnect_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( NastiRecursiveInterconnect_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( NastiRecursiveInterconnect_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( NastiRecursiveInterconnect_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( NastiRecursiveInterconnect_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( NastiRecursiveInterconnect_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( NastiRecursiveInterconnect_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( NastiRecursiveInterconnect_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( NastiRecursiveInterconnect_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( NastiRecursiveInterconnect_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( NastiRecursiveInterconnect_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( NastiRecursiveInterconnect_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( NastiRecursiveInterconnect_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( NastiRecursiveInterconnect_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( NastiRecursiveInterconnect_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( NastiRecursiveInterconnect_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( NastiRecursiveInterconnect_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiErrorSlave NastiErrorSlave(.clk(clk), .reset(reset),
       .io_aw_ready( NastiErrorSlave_io_aw_ready ),
       .io_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_w_ready( NastiErrorSlave_io_w_ready ),
       .io_w_valid( xbar_io_slaves_1_w_valid ),
       .io_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_b_ready( xbar_io_slaves_1_b_ready ),
       .io_b_valid( NastiErrorSlave_io_b_valid ),
       .io_b_bits_resp( NastiErrorSlave_io_b_bits_resp ),
       .io_b_bits_id( NastiErrorSlave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( NastiErrorSlave_io_ar_ready ),
       .io_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_r_ready( xbar_io_slaves_1_r_ready ),
       .io_r_valid( NastiErrorSlave_io_r_valid ),
       .io_r_bits_resp( NastiErrorSlave_io_r_bits_resp ),
       .io_r_bits_data( NastiErrorSlave_io_r_bits_data ),
       .io_r_bits_last( NastiErrorSlave_io_r_bits_last ),
       .io_r_bits_id( NastiErrorSlave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
endmodule

module NastiArbiter(
    output io_master_0_aw_ready,
    input  io_master_0_aw_valid,
    input [31:0] io_master_0_aw_bits_addr,
    input [7:0] io_master_0_aw_bits_len,
    input [2:0] io_master_0_aw_bits_size,
    input [1:0] io_master_0_aw_bits_burst,
    input  io_master_0_aw_bits_lock,
    input [3:0] io_master_0_aw_bits_cache,
    input [2:0] io_master_0_aw_bits_prot,
    input [3:0] io_master_0_aw_bits_qos,
    input [3:0] io_master_0_aw_bits_region,
    input [5:0] io_master_0_aw_bits_id,
    input  io_master_0_aw_bits_user,
    output io_master_0_w_ready,
    input  io_master_0_w_valid,
    input [63:0] io_master_0_w_bits_data,
    input  io_master_0_w_bits_last,
    input [7:0] io_master_0_w_bits_strb,
    input  io_master_0_w_bits_user,
    input  io_master_0_b_ready,
    output io_master_0_b_valid,
    output[1:0] io_master_0_b_bits_resp,
    output[5:0] io_master_0_b_bits_id,
    output io_master_0_b_bits_user,
    output io_master_0_ar_ready,
    input  io_master_0_ar_valid,
    input [31:0] io_master_0_ar_bits_addr,
    input [7:0] io_master_0_ar_bits_len,
    input [2:0] io_master_0_ar_bits_size,
    input [1:0] io_master_0_ar_bits_burst,
    input  io_master_0_ar_bits_lock,
    input [3:0] io_master_0_ar_bits_cache,
    input [2:0] io_master_0_ar_bits_prot,
    input [3:0] io_master_0_ar_bits_qos,
    input [3:0] io_master_0_ar_bits_region,
    input [5:0] io_master_0_ar_bits_id,
    input  io_master_0_ar_bits_user,
    input  io_master_0_r_ready,
    output io_master_0_r_valid,
    output[1:0] io_master_0_r_bits_resp,
    output[63:0] io_master_0_r_bits_data,
    output io_master_0_r_bits_last,
    output[5:0] io_master_0_r_bits_id,
    output io_master_0_r_bits_user,
    input  io_slave_aw_ready,
    output io_slave_aw_valid,
    output[31:0] io_slave_aw_bits_addr,
    output[7:0] io_slave_aw_bits_len,
    output[2:0] io_slave_aw_bits_size,
    output[1:0] io_slave_aw_bits_burst,
    output io_slave_aw_bits_lock,
    output[3:0] io_slave_aw_bits_cache,
    output[2:0] io_slave_aw_bits_prot,
    output[3:0] io_slave_aw_bits_qos,
    output[3:0] io_slave_aw_bits_region,
    output[5:0] io_slave_aw_bits_id,
    output io_slave_aw_bits_user,
    input  io_slave_w_ready,
    output io_slave_w_valid,
    output[63:0] io_slave_w_bits_data,
    output io_slave_w_bits_last,
    output[7:0] io_slave_w_bits_strb,
    output io_slave_w_bits_user,
    output io_slave_b_ready,
    input  io_slave_b_valid,
    input [1:0] io_slave_b_bits_resp,
    input [5:0] io_slave_b_bits_id,
    input  io_slave_b_bits_user,
    input  io_slave_ar_ready,
    output io_slave_ar_valid,
    output[31:0] io_slave_ar_bits_addr,
    output[7:0] io_slave_ar_bits_len,
    output[2:0] io_slave_ar_bits_size,
    output[1:0] io_slave_ar_bits_burst,
    output io_slave_ar_bits_lock,
    output[3:0] io_slave_ar_bits_cache,
    output[2:0] io_slave_ar_bits_prot,
    output[3:0] io_slave_ar_bits_qos,
    output[3:0] io_slave_ar_bits_region,
    output[5:0] io_slave_ar_bits_id,
    output io_slave_ar_bits_user,
    output io_slave_r_ready,
    input  io_slave_r_valid,
    input [1:0] io_slave_r_bits_resp,
    input [63:0] io_slave_r_bits_data,
    input  io_slave_r_bits_last,
    input [5:0] io_slave_r_bits_id,
    input  io_slave_r_bits_user
);



  assign io_slave_r_ready = io_master_0_r_ready;
  assign io_slave_ar_bits_user = io_master_0_ar_bits_user;
  assign io_slave_ar_bits_id = io_master_0_ar_bits_id;
  assign io_slave_ar_bits_region = io_master_0_ar_bits_region;
  assign io_slave_ar_bits_qos = io_master_0_ar_bits_qos;
  assign io_slave_ar_bits_prot = io_master_0_ar_bits_prot;
  assign io_slave_ar_bits_cache = io_master_0_ar_bits_cache;
  assign io_slave_ar_bits_lock = io_master_0_ar_bits_lock;
  assign io_slave_ar_bits_burst = io_master_0_ar_bits_burst;
  assign io_slave_ar_bits_size = io_master_0_ar_bits_size;
  assign io_slave_ar_bits_len = io_master_0_ar_bits_len;
  assign io_slave_ar_bits_addr = io_master_0_ar_bits_addr;
  assign io_slave_ar_valid = io_master_0_ar_valid;
  assign io_slave_b_ready = io_master_0_b_ready;
  assign io_slave_w_bits_user = io_master_0_w_bits_user;
  assign io_slave_w_bits_strb = io_master_0_w_bits_strb;
  assign io_slave_w_bits_last = io_master_0_w_bits_last;
  assign io_slave_w_bits_data = io_master_0_w_bits_data;
  assign io_slave_w_valid = io_master_0_w_valid;
  assign io_slave_aw_bits_user = io_master_0_aw_bits_user;
  assign io_slave_aw_bits_id = io_master_0_aw_bits_id;
  assign io_slave_aw_bits_region = io_master_0_aw_bits_region;
  assign io_slave_aw_bits_qos = io_master_0_aw_bits_qos;
  assign io_slave_aw_bits_prot = io_master_0_aw_bits_prot;
  assign io_slave_aw_bits_cache = io_master_0_aw_bits_cache;
  assign io_slave_aw_bits_lock = io_master_0_aw_bits_lock;
  assign io_slave_aw_bits_burst = io_master_0_aw_bits_burst;
  assign io_slave_aw_bits_size = io_master_0_aw_bits_size;
  assign io_slave_aw_bits_len = io_master_0_aw_bits_len;
  assign io_slave_aw_bits_addr = io_master_0_aw_bits_addr;
  assign io_slave_aw_valid = io_master_0_aw_valid;
  assign io_master_0_r_bits_user = io_slave_r_bits_user;
  assign io_master_0_r_bits_id = io_slave_r_bits_id;
  assign io_master_0_r_bits_last = io_slave_r_bits_last;
  assign io_master_0_r_bits_data = io_slave_r_bits_data;
  assign io_master_0_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_0_r_valid = io_slave_r_valid;
  assign io_master_0_ar_ready = io_slave_ar_ready;
  assign io_master_0_b_bits_user = io_slave_b_bits_user;
  assign io_master_0_b_bits_id = io_slave_b_bits_id;
  assign io_master_0_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_0_b_valid = io_slave_b_valid;
  assign io_master_0_w_ready = io_slave_w_ready;
  assign io_master_0_aw_ready = io_slave_aw_ready;
endmodule

module NastiMemoryInterconnect(
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [5:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[5:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [5:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[5:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[5:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [5:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[5:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [5:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiArbiter_io_master_0_aw_ready;
  wire NastiArbiter_io_master_0_w_ready;
  wire NastiArbiter_io_master_0_b_valid;
  wire[1:0] NastiArbiter_io_master_0_b_bits_resp;
  wire[5:0] NastiArbiter_io_master_0_b_bits_id;
  wire NastiArbiter_io_master_0_b_bits_user;
  wire NastiArbiter_io_master_0_ar_ready;
  wire NastiArbiter_io_master_0_r_valid;
  wire[1:0] NastiArbiter_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_0_r_bits_data;
  wire NastiArbiter_io_master_0_r_bits_last;
  wire[5:0] NastiArbiter_io_master_0_r_bits_id;
  wire NastiArbiter_io_master_0_r_bits_user;
  wire NastiArbiter_io_slave_aw_valid;
  wire[31:0] NastiArbiter_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_io_slave_aw_bits_burst;
  wire NastiArbiter_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_io_slave_aw_bits_region;
  wire[5:0] NastiArbiter_io_slave_aw_bits_id;
  wire NastiArbiter_io_slave_aw_bits_user;
  wire NastiArbiter_io_slave_w_valid;
  wire[63:0] NastiArbiter_io_slave_w_bits_data;
  wire NastiArbiter_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_io_slave_w_bits_strb;
  wire NastiArbiter_io_slave_w_bits_user;
  wire NastiArbiter_io_slave_b_ready;
  wire NastiArbiter_io_slave_ar_valid;
  wire[31:0] NastiArbiter_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_io_slave_ar_bits_burst;
  wire NastiArbiter_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_io_slave_ar_bits_region;
  wire[5:0] NastiArbiter_io_slave_ar_bits_id;
  wire NastiArbiter_io_slave_ar_bits_user;
  wire NastiArbiter_io_slave_r_ready;


  assign io_slaves_0_r_ready = NastiArbiter_io_slave_r_ready;
  assign io_slaves_0_ar_bits_user = NastiArbiter_io_slave_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiArbiter_io_slave_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiArbiter_io_slave_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiArbiter_io_slave_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiArbiter_io_slave_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiArbiter_io_slave_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiArbiter_io_slave_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiArbiter_io_slave_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiArbiter_io_slave_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiArbiter_io_slave_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiArbiter_io_slave_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiArbiter_io_slave_ar_valid;
  assign io_slaves_0_b_ready = NastiArbiter_io_slave_b_ready;
  assign io_slaves_0_w_bits_user = NastiArbiter_io_slave_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiArbiter_io_slave_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiArbiter_io_slave_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiArbiter_io_slave_w_bits_data;
  assign io_slaves_0_w_valid = NastiArbiter_io_slave_w_valid;
  assign io_slaves_0_aw_bits_user = NastiArbiter_io_slave_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiArbiter_io_slave_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiArbiter_io_slave_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiArbiter_io_slave_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiArbiter_io_slave_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiArbiter_io_slave_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiArbiter_io_slave_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiArbiter_io_slave_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiArbiter_io_slave_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiArbiter_io_slave_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiArbiter_io_slave_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiArbiter_io_slave_aw_valid;
  assign io_masters_0_r_bits_user = NastiArbiter_io_master_0_r_bits_user;
  assign io_masters_0_r_bits_id = NastiArbiter_io_master_0_r_bits_id;
  assign io_masters_0_r_bits_last = NastiArbiter_io_master_0_r_bits_last;
  assign io_masters_0_r_bits_data = NastiArbiter_io_master_0_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiArbiter_io_master_0_r_bits_resp;
  assign io_masters_0_r_valid = NastiArbiter_io_master_0_r_valid;
  assign io_masters_0_ar_ready = NastiArbiter_io_master_0_ar_ready;
  assign io_masters_0_b_bits_user = NastiArbiter_io_master_0_b_bits_user;
  assign io_masters_0_b_bits_id = NastiArbiter_io_master_0_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiArbiter_io_master_0_b_bits_resp;
  assign io_masters_0_b_valid = NastiArbiter_io_master_0_b_valid;
  assign io_masters_0_w_ready = NastiArbiter_io_master_0_w_ready;
  assign io_masters_0_aw_ready = NastiArbiter_io_master_0_aw_ready;
  NastiArbiter NastiArbiter(
       .io_master_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_master_0_aw_valid( io_masters_0_aw_valid ),
       .io_master_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_master_0_w_valid( io_masters_0_w_valid ),
       .io_master_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_0_b_ready( io_masters_0_b_ready ),
       .io_master_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_master_0_ar_valid( io_masters_0_ar_valid ),
       .io_master_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_0_r_ready( io_masters_0_r_ready ),
       .io_master_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_0_w_ready ),
       .io_slave_w_valid( NastiArbiter_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_0_b_valid ),
       .io_slave_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_0_r_valid ),
       .io_slave_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [3:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [3:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[3:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T54;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T55;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  locked;
  wire T56;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  reg [1:0] R20;
  wire[1:0] T57;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[127:0] T24;
  wire T25;
  wire[16:0] T26;
  wire[2:0] T27;
  wire T28;
  wire[1:0] T29;
  wire[3:0] T30;
  wire[25:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T54 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T55 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T14 & T12;
  assign T12 = io_out_bits_is_builtin_type & T13;
  assign T13 = 3'h3 == io_out_bits_a_type;
  assign T14 = io_out_valid & io_out_ready;
  assign T56 = reset ? 1'h0 : T15;
  assign T15 = T22 ? 1'h0 : T16;
  assign T16 = T11 ? T17 : locked;
  assign T17 = T18 ^ 1'h1;
  assign T18 = T19 == 2'h0;
  assign T19 = R20 + 2'h1;
  assign T57 = reset ? 2'h0 : T21;
  assign T21 = T11 ? T19 : R20;
  assign T22 = T14 & T23;
  assign T23 = T12 ^ 1'h1;
  assign io_out_bits_data = T24;
  assign T24 = T25 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T25 = chosen;
  assign io_out_bits_union = T26;
  assign T26 = T25 ? io_in_1_bits_union : io_in_0_bits_union;
  assign io_out_bits_a_type = T27;
  assign T27 = T25 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_is_builtin_type = T28;
  assign T28 = T25 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_addr_beat = T29;
  assign T29 = T25 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T30;
  assign T30 = T25 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T31;
  assign T31 = T25 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T32;
  assign T32 = T25 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T33;
  assign T33 = T34 & io_out_ready;
  assign T34 = locked ? T43 : T35;
  assign T35 = T42 | T36;
  assign T36 = T37 ^ 1'h1;
  assign T37 = T40 | T38;
  assign T38 = io_in_1_valid & T39;
  assign T39 = last_grant < 1'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = last_grant < 1'h0;
  assign T42 = last_grant < 1'h0;
  assign T43 = lockIdx == 1'h0;
  assign io_in_1_ready = T44;
  assign T44 = T45 & io_out_ready;
  assign T45 = locked ? T53 : T46;
  assign T46 = T50 | T47;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_0_valid;
  assign T49 = T40 | T38;
  assign T50 = T52 & T51;
  assign T51 = last_grant < 1'h1;
  assign T52 = T40 ^ 1'h1;
  assign T53 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T22) begin
      locked <= 1'h0;
    end else if(T11) begin
      locked <= T17;
    end
    if(reset) begin
      R20 <= 2'h0;
    end else if(T11) begin
      R20 <= T19;
    end
  end
endmodule

module ReorderQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_data,
    input [3:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [3:0] io_deq_tag,
    output io_deq_data,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_8;
  wire T1;
  reg  roq_free_8;
  wire T182;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[15:0] T6;
  wire[3:0] T7;
  wire[3:0] roq_enq_addr;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  reg  roq_free_7;
  wire T183;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[15:0] T21;
  wire[3:0] T22;
  wire[3:0] roq_deq_addr;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire roq_matches_7;
  wire T30;
  wire T31;
  reg [3:0] roq_tags_7;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire[15:0] T35;
  wire[3:0] T36;
  wire roq_matches_6;
  wire T37;
  wire T38;
  reg [3:0] roq_tags_6;
  wire[3:0] T39;
  wire T40;
  wire T41;
  wire roq_matches_5;
  wire T42;
  wire T43;
  reg [3:0] roq_tags_5;
  wire[3:0] T44;
  wire T45;
  wire T46;
  wire roq_matches_4;
  wire T47;
  wire T48;
  reg [3:0] roq_tags_4;
  wire[3:0] T49;
  wire T50;
  wire T51;
  wire roq_matches_3;
  wire T52;
  wire T53;
  reg [3:0] roq_tags_3;
  wire[3:0] T54;
  wire T55;
  wire T56;
  wire roq_matches_2;
  wire T57;
  wire T58;
  reg [3:0] roq_tags_2;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire roq_matches_1;
  wire T62;
  wire T63;
  reg [3:0] roq_tags_1;
  wire[3:0] T64;
  wire T65;
  wire T66;
  wire roq_matches_0;
  wire T67;
  wire T68;
  reg [3:0] roq_tags_0;
  wire[3:0] T69;
  wire T70;
  wire T71;
  reg  roq_free_6;
  wire T184;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  roq_free_5;
  wire T185;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  reg  roq_free_4;
  wire T186;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  roq_free_3;
  wire T187;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  roq_free_2;
  wire T188;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  reg  roq_free_1;
  wire T189;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  roq_free_0;
  wire T190;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  reg [3:0] roq_tags_8;
  wire[3:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg  roq_data_0;
  wire T132;
  wire T133;
  wire T134;
  wire[15:0] T135;
  wire[3:0] T136;
  reg  roq_data_1;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  reg  roq_data_2;
  wire T143;
  wire T144;
  wire T145;
  reg  roq_data_3;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  roq_data_4;
  wire T153;
  wire T154;
  wire T155;
  reg  roq_data_5;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  reg  roq_data_6;
  wire T161;
  wire T162;
  wire T163;
  reg  roq_data_7;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  reg  roq_data_8;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_8 = {1{$random}};
    roq_free_7 = {1{$random}};
    roq_tags_7 = {1{$random}};
    roq_tags_6 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_6 = {1{$random}};
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_8 = {1{$random}};
    roq_data_0 = {1{$random}};
    roq_data_1 = {1{$random}};
    roq_data_2 = {1{$random}};
    roq_data_3 = {1{$random}};
    roq_data_4 = {1{$random}};
    roq_data_5 = {1{$random}};
    roq_data_6 = {1{$random}};
    roq_data_7 = {1{$random}};
    roq_data_8 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T121 | roq_matches_8;
  assign roq_matches_8 = T117 & T1;
  assign T1 = roq_free_8 ^ 1'h1;
  assign T182 = reset ? 1'h1 : T2;
  assign T2 = T115 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_8;
  assign T4 = T114 & T5;
  assign T5 = T6[4'h8];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 4'h0 : T8;
  assign T8 = roq_free_1 ? 4'h1 : T9;
  assign T9 = roq_free_2 ? 4'h2 : T10;
  assign T10 = roq_free_3 ? 4'h3 : T11;
  assign T11 = roq_free_4 ? 4'h4 : T12;
  assign T12 = roq_free_5 ? 4'h5 : T13;
  assign T13 = roq_free_6 ? 4'h6 : T14;
  assign T14 = roq_free_7 ? 4'h7 : 4'h8;
  assign T183 = reset ? 1'h1 : T15;
  assign T15 = T19 ? 1'h1 : T16;
  assign T16 = T17 ? 1'h0 : roq_free_7;
  assign T17 = T114 & T18;
  assign T18 = T6[3'h7];
  assign T19 = io_deq_valid & T20;
  assign T20 = T21[3'h7];
  assign T21 = 1'h1 << T22;
  assign T22 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 4'h0 : T23;
  assign T23 = roq_matches_1 ? 4'h1 : T24;
  assign T24 = roq_matches_2 ? 4'h2 : T25;
  assign T25 = roq_matches_3 ? 4'h3 : T26;
  assign T26 = roq_matches_4 ? 4'h4 : T27;
  assign T27 = roq_matches_5 ? 4'h5 : T28;
  assign T28 = roq_matches_6 ? 4'h6 : T29;
  assign T29 = roq_matches_7 ? 4'h7 : 4'h8;
  assign roq_matches_7 = T31 & T30;
  assign T30 = roq_free_7 ^ 1'h1;
  assign T31 = roq_tags_7 == io_deq_tag;
  assign T32 = T33 ? io_enq_bits_tag : roq_tags_7;
  assign T33 = T114 & T34;
  assign T34 = T35[3'h7];
  assign T35 = 1'h1 << T36;
  assign T36 = roq_enq_addr;
  assign roq_matches_6 = T38 & T37;
  assign T37 = roq_free_6 ^ 1'h1;
  assign T38 = roq_tags_6 == io_deq_tag;
  assign T39 = T40 ? io_enq_bits_tag : roq_tags_6;
  assign T40 = T114 & T41;
  assign T41 = T35[3'h6];
  assign roq_matches_5 = T43 & T42;
  assign T42 = roq_free_5 ^ 1'h1;
  assign T43 = roq_tags_5 == io_deq_tag;
  assign T44 = T45 ? io_enq_bits_tag : roq_tags_5;
  assign T45 = T114 & T46;
  assign T46 = T35[3'h5];
  assign roq_matches_4 = T48 & T47;
  assign T47 = roq_free_4 ^ 1'h1;
  assign T48 = roq_tags_4 == io_deq_tag;
  assign T49 = T50 ? io_enq_bits_tag : roq_tags_4;
  assign T50 = T114 & T51;
  assign T51 = T35[3'h4];
  assign roq_matches_3 = T53 & T52;
  assign T52 = roq_free_3 ^ 1'h1;
  assign T53 = roq_tags_3 == io_deq_tag;
  assign T54 = T55 ? io_enq_bits_tag : roq_tags_3;
  assign T55 = T114 & T56;
  assign T56 = T35[2'h3];
  assign roq_matches_2 = T58 & T57;
  assign T57 = roq_free_2 ^ 1'h1;
  assign T58 = roq_tags_2 == io_deq_tag;
  assign T59 = T60 ? io_enq_bits_tag : roq_tags_2;
  assign T60 = T114 & T61;
  assign T61 = T35[2'h2];
  assign roq_matches_1 = T63 & T62;
  assign T62 = roq_free_1 ^ 1'h1;
  assign T63 = roq_tags_1 == io_deq_tag;
  assign T64 = T65 ? io_enq_bits_tag : roq_tags_1;
  assign T65 = T114 & T66;
  assign T66 = T35[1'h1];
  assign roq_matches_0 = T68 & T67;
  assign T67 = roq_free_0 ^ 1'h1;
  assign T68 = roq_tags_0 == io_deq_tag;
  assign T69 = T70 ? io_enq_bits_tag : roq_tags_0;
  assign T70 = T114 & T71;
  assign T71 = T35[1'h0];
  assign T184 = reset ? 1'h1 : T72;
  assign T72 = T76 ? 1'h1 : T73;
  assign T73 = T74 ? 1'h0 : roq_free_6;
  assign T74 = T114 & T75;
  assign T75 = T6[3'h6];
  assign T76 = io_deq_valid & T77;
  assign T77 = T21[3'h6];
  assign T185 = reset ? 1'h1 : T78;
  assign T78 = T82 ? 1'h1 : T79;
  assign T79 = T80 ? 1'h0 : roq_free_5;
  assign T80 = T114 & T81;
  assign T81 = T6[3'h5];
  assign T82 = io_deq_valid & T83;
  assign T83 = T21[3'h5];
  assign T186 = reset ? 1'h1 : T84;
  assign T84 = T88 ? 1'h1 : T85;
  assign T85 = T86 ? 1'h0 : roq_free_4;
  assign T86 = T114 & T87;
  assign T87 = T6[3'h4];
  assign T88 = io_deq_valid & T89;
  assign T89 = T21[3'h4];
  assign T187 = reset ? 1'h1 : T90;
  assign T90 = T94 ? 1'h1 : T91;
  assign T91 = T92 ? 1'h0 : roq_free_3;
  assign T92 = T114 & T93;
  assign T93 = T6[2'h3];
  assign T94 = io_deq_valid & T95;
  assign T95 = T21[2'h3];
  assign T188 = reset ? 1'h1 : T96;
  assign T96 = T100 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : roq_free_2;
  assign T98 = T114 & T99;
  assign T99 = T6[2'h2];
  assign T100 = io_deq_valid & T101;
  assign T101 = T21[2'h2];
  assign T189 = reset ? 1'h1 : T102;
  assign T102 = T106 ? 1'h1 : T103;
  assign T103 = T104 ? 1'h0 : roq_free_1;
  assign T104 = T114 & T105;
  assign T105 = T6[1'h1];
  assign T106 = io_deq_valid & T107;
  assign T107 = T21[1'h1];
  assign T190 = reset ? 1'h1 : T108;
  assign T108 = T112 ? 1'h1 : T109;
  assign T109 = T110 ? 1'h0 : roq_free_0;
  assign T110 = T114 & T111;
  assign T111 = T6[1'h0];
  assign T112 = io_deq_valid & T113;
  assign T113 = T21[1'h0];
  assign T114 = io_enq_valid & io_enq_ready;
  assign T115 = io_deq_valid & T116;
  assign T116 = T21[4'h8];
  assign T117 = roq_tags_8 == io_deq_tag;
  assign T118 = T119 ? io_enq_bits_tag : roq_tags_8;
  assign T119 = T114 & T120;
  assign T120 = T35[4'h8];
  assign T121 = T122 | roq_matches_7;
  assign T122 = T123 | roq_matches_6;
  assign T123 = T124 | roq_matches_5;
  assign T124 = T125 | roq_matches_4;
  assign T125 = T126 | roq_matches_3;
  assign T126 = T127 | roq_matches_2;
  assign T127 = roq_matches_0 | roq_matches_1;
  assign io_deq_data = T128;
  assign T128 = T173 ? roq_data_8 : T129;
  assign T129 = T169 ? T151 : T130;
  assign T130 = T150 ? T142 : T131;
  assign T131 = T140 ? roq_data_1 : roq_data_0;
  assign T132 = T133 ? io_enq_bits_data : roq_data_0;
  assign T133 = T114 & T134;
  assign T134 = T135[1'h0];
  assign T135 = 1'h1 << T136;
  assign T136 = roq_enq_addr;
  assign T137 = T138 ? io_enq_bits_data : roq_data_1;
  assign T138 = T114 & T139;
  assign T139 = T135[1'h1];
  assign T140 = T141[1'h0];
  assign T141 = roq_deq_addr;
  assign T142 = T149 ? roq_data_3 : roq_data_2;
  assign T143 = T144 ? io_enq_bits_data : roq_data_2;
  assign T144 = T114 & T145;
  assign T145 = T135[2'h2];
  assign T146 = T147 ? io_enq_bits_data : roq_data_3;
  assign T147 = T114 & T148;
  assign T148 = T135[2'h3];
  assign T149 = T141[1'h0];
  assign T150 = T141[1'h1];
  assign T151 = T168 ? T160 : T152;
  assign T152 = T159 ? roq_data_5 : roq_data_4;
  assign T153 = T154 ? io_enq_bits_data : roq_data_4;
  assign T154 = T114 & T155;
  assign T155 = T135[3'h4];
  assign T156 = T157 ? io_enq_bits_data : roq_data_5;
  assign T157 = T114 & T158;
  assign T158 = T135[3'h5];
  assign T159 = T141[1'h0];
  assign T160 = T167 ? roq_data_7 : roq_data_6;
  assign T161 = T162 ? io_enq_bits_data : roq_data_6;
  assign T162 = T114 & T163;
  assign T163 = T135[3'h6];
  assign T164 = T165 ? io_enq_bits_data : roq_data_7;
  assign T165 = T114 & T166;
  assign T166 = T135[3'h7];
  assign T167 = T141[1'h0];
  assign T168 = T141[1'h1];
  assign T169 = T141[2'h2];
  assign T170 = T171 ? io_enq_bits_data : roq_data_8;
  assign T171 = T114 & T172;
  assign T172 = T135[4'h8];
  assign T173 = T141[2'h3];
  assign io_enq_ready = T174;
  assign T174 = T175 | roq_free_8;
  assign T175 = T176 | roq_free_7;
  assign T176 = T177 | roq_free_6;
  assign T177 = T178 | roq_free_5;
  assign T178 = T179 | roq_free_4;
  assign T179 = T180 | roq_free_3;
  assign T180 = T181 | roq_free_2;
  assign T181 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_8 <= 1'h1;
    end else if(T115) begin
      roq_free_8 <= 1'h1;
    end else if(T4) begin
      roq_free_8 <= 1'h0;
    end
    if(reset) begin
      roq_free_7 <= 1'h1;
    end else if(T19) begin
      roq_free_7 <= 1'h1;
    end else if(T17) begin
      roq_free_7 <= 1'h0;
    end
    if(T33) begin
      roq_tags_7 <= io_enq_bits_tag;
    end
    if(T40) begin
      roq_tags_6 <= io_enq_bits_tag;
    end
    if(T45) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T50) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T55) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T60) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T65) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T70) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_6 <= 1'h1;
    end else if(T76) begin
      roq_free_6 <= 1'h1;
    end else if(T74) begin
      roq_free_6 <= 1'h0;
    end
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T82) begin
      roq_free_5 <= 1'h1;
    end else if(T80) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T88) begin
      roq_free_4 <= 1'h1;
    end else if(T86) begin
      roq_free_4 <= 1'h0;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T94) begin
      roq_free_3 <= 1'h1;
    end else if(T92) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T100) begin
      roq_free_2 <= 1'h1;
    end else if(T98) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T106) begin
      roq_free_1 <= 1'h1;
    end else if(T104) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T112) begin
      roq_free_0 <= 1'h1;
    end else if(T110) begin
      roq_free_0 <= 1'h0;
    end
    if(T119) begin
      roq_tags_8 <= io_enq_bits_tag;
    end
    if(T133) begin
      roq_data_0 <= io_enq_bits_data;
    end
    if(T138) begin
      roq_data_1 <= io_enq_bits_data;
    end
    if(T144) begin
      roq_data_2 <= io_enq_bits_data;
    end
    if(T147) begin
      roq_data_3 <= io_enq_bits_data;
    end
    if(T154) begin
      roq_data_4 <= io_enq_bits_data;
    end
    if(T157) begin
      roq_data_5 <= io_enq_bits_data;
    end
    if(T162) begin
      roq_data_6 <= io_enq_bits_data;
    end
    if(T165) begin
      roq_data_7 <= io_enq_bits_data;
    end
    if(T171) begin
      roq_data_8 <= io_enq_bits_data;
    end
  end
endmodule

module ClientTileLinkIOUnwrapper(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_in_probe_ready,
    output io_in_probe_valid,
    //output[25:0] io_in_probe_bits_addr_block
    //output[1:0] io_in_probe_bits_p_type
    output io_in_release_ready,
    input  io_in_release_valid,
    input [1:0] io_in_release_bits_addr_beat,
    input [25:0] io_in_release_bits_addr_block,
    input [3:0] io_in_release_bits_client_xact_id,
    input  io_in_release_bits_voluntary,
    input [2:0] io_in_release_bits_r_type,
    input [127:0] io_in_release_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire rel_roq_enq;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire acq_roq_enq;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[127:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire T36;
  wire[1:0] T37;
  wire[3:0] T38;
  wire[25:0] T39;
  wire T40;
  wire acq_roq_ready;
  wire T41;
  wire[127:0] T42;
  wire[16:0] T43;
  wire[16:0] T44;
  wire[15:0] T45;
  wire[2:0] T46;
  wire T47;
  wire[1:0] T48;
  wire[3:0] T49;
  wire[25:0] T50;
  wire T51;
  wire rel_roq_ready;
  wire T52;
  wire T53;
  wire[127:0] T54;
  wire[127:0] rel_grant_data;
  wire[127:0] acq_grant_data;
  wire[3:0] T55;
  wire[3:0] rel_grant_g_type;
  wire[3:0] T56;
  wire[3:0] acq_grant_g_type;
  wire[3:0] T57;
  wire T58;
  wire rel_grant_is_builtin_type;
  wire acq_grant_is_builtin_type;
  wire T59;
  wire rel_grant_manager_xact_id;
  wire acq_grant_manager_xact_id;
  wire[3:0] T60;
  wire[3:0] rel_grant_client_xact_id;
  wire[3:0] acq_grant_client_xact_id;
  wire[1:0] T61;
  wire[1:0] rel_grant_addr_beat;
  wire[1:0] acq_grant_addr_beat;
  wire T62;
  wire acqArb_io_in_1_ready;
  wire acqArb_io_in_0_ready;
  wire acqArb_io_out_valid;
  wire[25:0] acqArb_io_out_bits_addr_block;
  wire[3:0] acqArb_io_out_bits_client_xact_id;
  wire[1:0] acqArb_io_out_bits_addr_beat;
  wire acqArb_io_out_bits_is_builtin_type;
  wire[2:0] acqArb_io_out_bits_a_type;
  wire[16:0] acqArb_io_out_bits_union;
  wire[127:0] acqArb_io_out_bits_data;
  wire acqRoq_io_enq_ready;
  wire acqRoq_io_deq_data;
  wire acqRoq_io_deq_matches;
  wire relRoq_io_enq_ready;
  wire relRoq_io_deq_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_in_probe_bits_p_type = {1{$random}};
//  assign io_in_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T7 & T1;
  assign T1 = T3 | T2;
  assign T2 = io_out_grant_bits_addr_beat == 2'h3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = io_out_grant_bits_is_builtin_type ? T6 : T5;
  assign T5 = 4'h0 == io_out_grant_bits_g_type;
  assign T6 = 4'h5 == io_out_grant_bits_g_type;
  assign T7 = io_out_grant_ready & io_out_grant_valid;
  assign T8 = T16 & rel_roq_enq;
  assign rel_roq_enq = T10 | T9;
  assign T9 = io_in_release_bits_addr_beat == 2'h0;
  assign T10 = T11 ^ 1'h1;
  assign T11 = T13 | T12;
  assign T12 = 3'h2 == io_in_release_bits_r_type;
  assign T13 = T15 | T14;
  assign T14 = 3'h1 == io_in_release_bits_r_type;
  assign T15 = 3'h0 == io_in_release_bits_r_type;
  assign T16 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T17 = T24 & T18;
  assign T18 = T20 | T19;
  assign T19 = io_out_grant_bits_addr_beat == 2'h3;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_out_grant_bits_is_builtin_type ? T23 : T22;
  assign T22 = 4'h0 == io_out_grant_bits_g_type;
  assign T23 = 4'h5 == io_out_grant_bits_g_type;
  assign T24 = io_out_grant_ready & io_out_grant_valid;
  assign T25 = T30 & acq_roq_enq;
  assign acq_roq_enq = T27 | T26;
  assign T26 = io_in_acquire_bits_addr_beat == 2'h0;
  assign T27 = T28 ^ 1'h1;
  assign T28 = io_in_acquire_bits_is_builtin_type & T29;
  assign T29 = 3'h3 == io_in_acquire_bits_a_type;
  assign T30 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T31 = io_in_acquire_bits_data;
  assign T32 = T33;
  assign T33 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : 17'h1c1;
  assign T34 = T35;
  assign T35 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T36 = 1'h1;
  assign T37 = io_in_acquire_bits_addr_beat;
  assign T38 = io_in_acquire_bits_client_xact_id;
  assign T39 = io_in_acquire_bits_addr_block;
  assign T40 = io_in_acquire_valid & acq_roq_ready;
  assign acq_roq_ready = T41 | acqRoq_io_enq_ready;
  assign T41 = acq_roq_enq ^ 1'h1;
  assign T42 = io_in_release_bits_data;
  assign T43 = T44;
  assign T44 = {T45, 1'h1};
  assign T45 = 16'hffff;
  assign T46 = 3'h3;
  assign T47 = 1'h1;
  assign T48 = io_in_release_bits_addr_beat;
  assign T49 = io_in_release_bits_client_xact_id;
  assign T50 = io_in_release_bits_addr_block;
  assign T51 = io_in_release_valid & rel_roq_ready;
  assign rel_roq_ready = T52 | relRoq_io_enq_ready;
  assign T52 = rel_roq_enq ^ 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_in_release_ready = T53;
  assign T53 = rel_roq_ready & acqArb_io_in_1_ready;
  assign io_in_probe_valid = 1'h0;
  assign io_in_grant_bits_data = T54;
  assign T54 = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
  assign rel_grant_data = io_out_grant_bits_data;
  assign acq_grant_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = T55;
  assign T55 = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign rel_grant_g_type = T56;
  assign T56 = relRoq_io_deq_data ? 4'h0 : io_out_grant_bits_g_type;
  assign acq_grant_g_type = T57;
  assign T57 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign io_in_grant_bits_is_builtin_type = T58;
  assign T58 = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign rel_grant_is_builtin_type = 1'h1;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign io_in_grant_bits_manager_xact_id = T59;
  assign T59 = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = T60;
  assign T60 = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = T61;
  assign T61 = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = T62;
  assign T62 = acq_roq_ready & acqArb_io_in_0_ready;
  LockingRRArbiter_4 acqArb(.clk(clk), .reset(reset),
       .io_in_1_ready( acqArb_io_in_1_ready ),
       .io_in_1_valid( T51 ),
       .io_in_1_bits_addr_block( T50 ),
       .io_in_1_bits_client_xact_id( T49 ),
       .io_in_1_bits_addr_beat( T48 ),
       .io_in_1_bits_is_builtin_type( T47 ),
       .io_in_1_bits_a_type( T46 ),
       .io_in_1_bits_union( T43 ),
       .io_in_1_bits_data( T42 ),
       .io_in_0_ready( acqArb_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_addr_block( T39 ),
       .io_in_0_bits_client_xact_id( T38 ),
       .io_in_0_bits_addr_beat( T37 ),
       .io_in_0_bits_is_builtin_type( T36 ),
       .io_in_0_bits_a_type( T34 ),
       .io_in_0_bits_union( T32 ),
       .io_in_0_bits_data( T31 ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( acqArb_io_out_valid ),
       .io_out_bits_addr_block( acqArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( acqArb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( acqArb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( acqArb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( acqArb_io_out_bits_a_type ),
       .io_out_bits_union( acqArb_io_out_bits_union ),
       .io_out_bits_data( acqArb_io_out_bits_data )
       //.io_chosen(  )
  );
  ReorderQueue_0 acqRoq(.clk(clk), .reset(reset),
       .io_enq_ready( acqRoq_io_enq_ready ),
       .io_enq_valid( T25 ),
       .io_enq_bits_data( io_in_acquire_bits_is_builtin_type ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T17 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( acqRoq_io_deq_data ),
       .io_deq_matches( acqRoq_io_deq_matches )
  );
  ReorderQueue_0 relRoq(.clk(clk), .reset(reset),
       .io_enq_ready( relRoq_io_enq_ready ),
       .io_enq_valid( T8 ),
       .io_enq_bits_data( io_in_release_bits_voluntary ),
       .io_enq_bits_tag( io_in_release_bits_client_xact_id ),
       .io_deq_valid( T0 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( relRoq_io_deq_data )
       //.io_deq_matches(  )
  );
endmodule

module TileLinkIONarrower(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[2:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[11:0] io_out_acquire_bits_union,
    output[63:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [2:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [63:0] io_out_grant_bits_data
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire[1:0] T28;
  wire T29;
  wire[7:0] T30;
  wire[15:0] T31;
  wire[15:0] T32;
  wire[15:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[15:0] T39;
  wire[15:0] T40;
  wire[7:0] T41;
  wire[7:0] T318;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[3:0] T45;
  wire[7:0] T46;
  wire[7:0] T319;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[7:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[15:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire[15:0] T60;
  wire[15:0] T61;
  wire[7:0] T62;
  wire[7:0] T320;
  wire T63;
  wire[1:0] T64;
  wire T65;
  wire[3:0] T66;
  wire[7:0] T67;
  wire[7:0] T321;
  wire T68;
  wire T69;
  wire T70;
  wire[1:0] T322;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[31:0] T80;
  wire[5:0] T81;
  wire[3:0] T82;
  wire T83;
  wire T84;
  reg  R85;
  wire T323;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg  R93;
  wire T324;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg  R105;
  wire T325;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg  R110;
  wire T326;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[63:0] T327;
  wire[127:0] T117;
  wire[127:0] T118;
  wire[127:0] T119;
  wire[127:0] T120;
  wire[127:0] T121;
  wire[127:0] T328;
  wire[63:0] T122;
  wire[127:0] T329;
  wire[63:0] T123;
  wire[63:0] T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire[63:0] T128;
  wire[63:0] T129;
  wire T130;
  wire[127:0] T330;
  wire[63:0] T131;
  wire T132;
  wire[127:0] T331;
  wire[63:0] T133;
  wire[63:0] T134;
  reg [127:0] R135;
  wire[127:0] T136;
  wire[127:0] T137;
  wire[127:0] T332;
  wire[63:0] T138;
  wire[11:0] T333;
  wire[16:0] T139;
  wire[16:0] T140;
  wire[16:0] T141;
  wire[16:0] T142;
  wire[16:0] T143;
  wire[16:0] T334;
  wire[11:0] T144;
  wire[11:0] T145;
  wire[5:0] T146;
  wire T147;
  wire[5:0] T148;
  wire[2:0] T149;
  wire[2:0] T150;
  wire[31:0] T151;
  wire[5:0] T152;
  wire[3:0] T153;
  wire[16:0] T335;
  wire[11:0] T154;
  wire[11:0] T336;
  wire[8:0] T155;
  wire[7:0] T156;
  wire[7:0] T157;
  wire T158;
  wire[7:0] T159;
  wire T160;
  wire[16:0] T337;
  wire[11:0] T161;
  wire[11:0] T338;
  wire[8:0] T162;
  wire[5:0] T163;
  wire T164;
  wire[16:0] T339;
  wire[11:0] T165;
  wire[11:0] T340;
  wire[8:0] T166;
  wire[7:0] T167;
  reg [15:0] R168;
  wire[15:0] T169;
  wire[15:0] T170;
  wire[15:0] T171;
  wire[15:0] T172;
  wire[15:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire[15:0] T179;
  wire[15:0] T180;
  wire[7:0] T181;
  wire[7:0] T341;
  wire T182;
  wire[1:0] T183;
  wire T184;
  wire[3:0] T185;
  wire[7:0] T186;
  wire[7:0] T342;
  wire T187;
  wire T188;
  wire T189;
  wire[15:0] T343;
  wire[7:0] T190;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[2:0] T196;
  wire[2:0] T197;
  wire[2:0] T198;
  wire[2:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire[2:0] T209;
  wire[2:0] T210;
  wire[2:0] T211;
  wire[2:0] T212;
  wire[2:0] T344;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire[31:0] T216;
  wire[5:0] T217;
  wire[3:0] T218;
  wire[2:0] T219;
  wire[2:0] T220;
  wire T345;
  wire T346;
  wire[2:0] T222;
  wire[2:0] T223;
  wire[2:0] T224;
  reg [1:0] R225;
  wire[1:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[3:0] T230;
  wire[3:0] T231;
  wire[3:0] T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  reg [3:0] R236;
  wire[3:0] T237;
  wire[25:0] T238;
  wire[25:0] T239;
  wire[25:0] T240;
  wire[25:0] T241;
  wire[25:0] T242;
  wire[25:0] T243;
  wire[25:0] T244;
  wire[25:0] T245;
  wire[25:0] T246;
  reg [25:0] R247;
  wire[25:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[127:0] T256;
  wire[127:0] T257;
  wire[127:0] T347;
  wire[63:0] T258;
  wire[127:0] T259;
  wire[127:0] T348;
  wire[190:0] T260;
  wire[6:0] T261;
  wire[127:0] T262;
  wire[127:0] T263;
  wire[127:0] T264;
  reg [63:0] R265;
  wire[63:0] T266;
  wire T267;
  wire T268;
  wire[1:0] T269;
  wire T270;
  reg [63:0] R271;
  wire[63:0] T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[3:0] T278;
  wire[3:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  reg  R290;
  wire T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[3:0] T296;
  reg [3:0] R297;
  wire[3:0] T298;
  wire[1:0] T349;
  wire[2:0] T299;
  wire[2:0] T300;
  wire[2:0] T301;
  wire[2:0] T350;
  wire[1:0] T302;
  wire[1:0] T303;
  wire[2:0] T351;
  wire[1:0] T304;
  reg [1:0] R305;
  wire[1:0] T352;
  wire[1:0] T306;
  wire[1:0] T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire ReorderQueue_io_enq_ready;
  wire ReorderQueue_io_deq_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T21 = 1'b0;
    R85 = {1{$random}};
    R93 = {1{$random}};
    R105 = {1{$random}};
    R110 = {1{$random}};
    R135 = {4{$random}};
    R168 = {1{$random}};
    R225 = {1{$random}};
    R236 = {1{$random}};
    R247 = {1{$random}};
    R265 = {2{$random}};
    R271 = {2{$random}};
    R290 = {1{$random}};
    R297 = {1{$random}};
    R305 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T17 | T3;
  assign T3 = T16 ? 1'h1 : T4;
  assign T4 = T15 ? 1'h1 : T5;
  assign T5 = T14 ? 1'h1 : T6;
  assign T6 = T13 ? 1'h1 : T7;
  assign T7 = T12 ? 1'h1 : T8;
  assign T8 = T11 ? 1'h1 : T9;
  assign T9 = T10 == 3'h3;
  assign T10 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T11 = T10 == 3'h6;
  assign T12 = T10 == 3'h2;
  assign T13 = T10 == 3'h5;
  assign T14 = T10 == 3'h1;
  assign T15 = T10 == 3'h4;
  assign T16 = T10 == 3'h0;
  assign T17 = T20 | T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = io_in_acquire_bits_a_type == 3'h0;
  assign T20 = io_in_acquire_valid ^ 1'h1;
  assign T22 = T23 | reset;
  assign T23 = T72 | T24;
  assign T24 = T25 <= 2'h1;
  assign T25 = T322 + T26;
  assign T26 = {1'h0, T27};
  assign T27 = T28[1'h1];
  assign T28 = {T50, T29};
  assign T29 = T30 != 8'h0;
  assign T30 = T31[3'h7:1'h0];
  assign T31 = T48 ? T39 : T32;
  assign T32 = T34 ? T33 : 16'h0;
  assign T33 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T34 = T37 | T35;
  assign T35 = io_in_acquire_bits_is_builtin_type & T36;
  assign T36 = io_in_acquire_bits_a_type == 3'h2;
  assign T37 = io_in_acquire_bits_is_builtin_type & T38;
  assign T38 = io_in_acquire_bits_a_type == 3'h3;
  assign T39 = T40;
  assign T40 = {T46, T41};
  assign T41 = 8'h0 - T318;
  assign T318 = {7'h0, T42};
  assign T42 = T43[1'h0];
  assign T43 = 1'h1 << T44;
  assign T44 = T45[2'h3];
  assign T45 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T46 = 8'h0 - T319;
  assign T319 = {7'h0, T47};
  assign T47 = T43[1'h1];
  assign T48 = io_in_acquire_bits_is_builtin_type & T49;
  assign T49 = io_in_acquire_bits_a_type == 3'h4;
  assign T50 = T51 != 8'h0;
  assign T51 = T52[4'hf:4'h8];
  assign T52 = T69 ? T60 : T53;
  assign T53 = T55 ? T54 : 16'h0;
  assign T54 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T55 = T58 | T56;
  assign T56 = io_in_acquire_bits_is_builtin_type & T57;
  assign T57 = io_in_acquire_bits_a_type == 3'h2;
  assign T58 = io_in_acquire_bits_is_builtin_type & T59;
  assign T59 = io_in_acquire_bits_a_type == 3'h3;
  assign T60 = T61;
  assign T61 = {T67, T62};
  assign T62 = 8'h0 - T320;
  assign T320 = {7'h0, T63};
  assign T63 = T64[1'h0];
  assign T64 = 1'h1 << T65;
  assign T65 = T66[2'h3];
  assign T66 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T67 = 8'h0 - T321;
  assign T321 = {7'h0, T68};
  assign T68 = T64[1'h1];
  assign T69 = io_in_acquire_bits_is_builtin_type & T70;
  assign T70 = io_in_acquire_bits_a_type == 3'h4;
  assign T322 = {1'h0, T71};
  assign T71 = T28[1'h0];
  assign T72 = T75 | T73;
  assign T73 = T74 ^ 1'h1;
  assign T74 = io_in_acquire_bits_a_type == 3'h2;
  assign T75 = io_in_acquire_valid ^ 1'h1;
  assign T76 = T78 & T77;
  assign T77 = io_out_grant_bits_g_type == 4'h4;
  assign T78 = io_out_grant_ready & io_out_grant_valid;
  assign T79 = T80[2'h3];
  assign T80 = {io_in_acquire_bits_addr_block, T81};
  assign T81 = {io_in_acquire_bits_addr_beat, T82};
  assign T82 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T83 = T97 & T84;
  assign T84 = R85 ^ 1'h1;
  assign T323 = reset ? 1'h0 : T86;
  assign T86 = T91 ? 1'h0 : T87;
  assign T87 = T88 ? 1'h1 : R85;
  assign T88 = T90 & T89;
  assign T89 = io_in_acquire_bits_a_type == 3'h3;
  assign T90 = io_in_acquire_ready & io_in_acquire_valid;
  assign T91 = T96 & T92;
  assign T92 = R93 == 1'h1;
  assign T324 = reset ? 1'h0 : T94;
  assign T94 = T96 ? T95 : R93;
  assign T95 = R93 + 1'h1;
  assign T96 = R85 & io_out_acquire_ready;
  assign T97 = T98 & io_out_acquire_ready;
  assign T98 = T19 & io_in_acquire_valid;
  assign io_out_grant_ready = T99;
  assign T99 = T104 & T100;
  assign T100 = T101 | io_in_grant_ready;
  assign T101 = io_out_grant_bits_is_builtin_type ? T103 : T102;
  assign T102 = 4'h0 == io_out_grant_bits_g_type;
  assign T103 = 4'h5 == io_out_grant_bits_g_type;
  assign T104 = R105 ^ 1'h1;
  assign T325 = reset ? 1'h0 : T106;
  assign T106 = T116 ? 1'h0 : T107;
  assign T107 = T108 ? 1'h1 : R105;
  assign T108 = T113 & T109;
  assign T109 = R110 == 1'h1;
  assign T326 = reset ? 1'h0 : T111;
  assign T111 = T113 ? T112 : R110;
  assign T112 = R110 + 1'h1;
  assign T113 = T115 & T114;
  assign T114 = R105 ^ 1'h1;
  assign T115 = io_out_grant_valid & T101;
  assign T116 = io_in_grant_ready & R105;
  assign io_out_acquire_bits_data = T327;
  assign T327 = T117[6'h3f:1'h0];
  assign T117 = R85 ? T331 : T118;
  assign T118 = T132 ? T330 : T119;
  assign T119 = T74 ? T329 : T120;
  assign T120 = T19 ? T328 : T121;
  assign T121 = io_in_acquire_bits_data;
  assign T328 = {64'h0, T122};
  assign T122 = 64'h0;
  assign T329 = {64'h0, T123};
  assign T123 = T124;
  assign T124 = T128 | T125;
  assign T125 = T127 ? T126 : 64'h0;
  assign T126 = io_in_acquire_bits_data[7'h7f:7'h40];
  assign T127 = T28[1'h1];
  assign T128 = T130 ? T129 : 64'h0;
  assign T129 = io_in_acquire_bits_data[6'h3f:1'h0];
  assign T130 = T28[1'h0];
  assign T330 = {64'h0, T131};
  assign T131 = 64'h0;
  assign T132 = io_in_acquire_bits_a_type == 3'h1;
  assign T331 = {64'h0, T133};
  assign T133 = T134;
  assign T134 = R135[6'h3f:1'h0];
  assign T136 = T96 ? T332 : T137;
  assign T137 = T88 ? io_in_acquire_bits_data : R135;
  assign T332 = {64'h0, T138};
  assign T138 = R135 >> 7'h40;
  assign io_out_acquire_bits_union = T333;
  assign T333 = T139[4'hb:1'h0];
  assign T139 = R85 ? T339 : T140;
  assign T140 = T132 ? T337 : T141;
  assign T141 = T74 ? T335 : T142;
  assign T142 = T19 ? T334 : T143;
  assign T143 = io_in_acquire_bits_union;
  assign T334 = {5'h0, T144};
  assign T144 = T145;
  assign T145 = {T148, T146};
  assign T146 = {5'h0, T147};
  assign T147 = io_in_acquire_bits_union[1'h0];
  assign T148 = {T150, T149};
  assign T149 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T150 = T151[2'h2:1'h0];
  assign T151 = {io_in_acquire_bits_addr_block, T152};
  assign T152 = {io_in_acquire_bits_addr_beat, T153};
  assign T153 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T335 = {5'h0, T154};
  assign T154 = T336;
  assign T336 = {3'h0, T155};
  assign T155 = {T156, 1'h1};
  assign T156 = T159 | T157;
  assign T157 = T158 ? T51 : 8'h0;
  assign T158 = T28[1'h1];
  assign T159 = T160 ? T30 : 8'h0;
  assign T160 = T28[1'h0];
  assign T337 = {5'h0, T161};
  assign T161 = T338;
  assign T338 = {3'h0, T162};
  assign T162 = {3'h7, T163};
  assign T163 = {5'h0, T164};
  assign T164 = io_in_acquire_bits_union[1'h0];
  assign T339 = {5'h0, T165};
  assign T165 = T340;
  assign T340 = {3'h0, T166};
  assign T166 = {T167, 1'h1};
  assign T167 = R168[3'h7:1'h0];
  assign T169 = T96 ? T343 : T170;
  assign T170 = T88 ? T171 : R168;
  assign T171 = T188 ? T179 : T172;
  assign T172 = T174 ? T173 : 16'h0;
  assign T173 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T174 = T177 | T175;
  assign T175 = io_in_acquire_bits_is_builtin_type & T176;
  assign T176 = io_in_acquire_bits_a_type == 3'h2;
  assign T177 = io_in_acquire_bits_is_builtin_type & T178;
  assign T178 = io_in_acquire_bits_a_type == 3'h3;
  assign T179 = T180;
  assign T180 = {T186, T181};
  assign T181 = 8'h0 - T341;
  assign T341 = {7'h0, T182};
  assign T182 = T183[1'h0];
  assign T183 = 1'h1 << T184;
  assign T184 = T185[2'h3];
  assign T185 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T186 = 8'h0 - T342;
  assign T342 = {7'h0, T187};
  assign T187 = T183[1'h1];
  assign T188 = io_in_acquire_bits_is_builtin_type & T189;
  assign T189 = io_in_acquire_bits_a_type == 3'h4;
  assign T343 = {8'h0, T190};
  assign T190 = R168 >> 4'h8;
  assign io_out_acquire_bits_a_type = T191;
  assign T191 = R85 ? T199 : T192;
  assign T192 = T132 ? T198 : T193;
  assign T193 = T74 ? T197 : T194;
  assign T194 = T19 ? T196 : T195;
  assign T195 = io_in_acquire_bits_a_type;
  assign T196 = 3'h0;
  assign T197 = 3'h2;
  assign T198 = 3'h1;
  assign T199 = 3'h3;
  assign io_out_acquire_bits_is_builtin_type = T200;
  assign T200 = R85 ? T208 : T201;
  assign T201 = T132 ? T207 : T202;
  assign T202 = T74 ? T206 : T203;
  assign T203 = T19 ? T205 : T204;
  assign T204 = io_in_acquire_bits_is_builtin_type;
  assign T205 = 1'h1;
  assign T206 = 1'h1;
  assign T207 = 1'h1;
  assign T208 = 1'h1;
  assign io_out_acquire_bits_addr_beat = T209;
  assign T209 = R85 ? T223 : T210;
  assign T210 = T132 ? T222 : T211;
  assign T211 = T74 ? T219 : T212;
  assign T212 = T19 ? T214 : T344;
  assign T344 = {1'h0, T213};
  assign T213 = io_in_acquire_bits_addr_beat;
  assign T214 = T215;
  assign T215 = T216[3'h5:2'h3];
  assign T216 = {io_in_acquire_bits_addr_block, T217};
  assign T217 = {io_in_acquire_bits_addr_beat, T218};
  assign T218 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T219 = T220;
  assign T220 = {io_in_acquire_bits_addr_beat, T345};
  assign T345 = T346 == 1'h0;
  assign T346 = T28[1'h0];
  assign T222 = 3'h0;
  assign T223 = T224;
  assign T224 = {R225, R93};
  assign T226 = T88 ? io_in_acquire_bits_addr_beat : R225;
  assign io_out_acquire_bits_client_xact_id = T227;
  assign T227 = R85 ? T235 : T228;
  assign T228 = T132 ? T234 : T229;
  assign T229 = T74 ? T233 : T230;
  assign T230 = T19 ? T232 : T231;
  assign T231 = io_in_acquire_bits_client_xact_id;
  assign T232 = io_in_acquire_bits_client_xact_id;
  assign T233 = io_in_acquire_bits_client_xact_id;
  assign T234 = io_in_acquire_bits_client_xact_id;
  assign T235 = R236;
  assign T237 = T88 ? io_in_acquire_bits_client_xact_id : R236;
  assign io_out_acquire_bits_addr_block = T238;
  assign T238 = R85 ? T246 : T239;
  assign T239 = T132 ? T245 : T240;
  assign T240 = T74 ? T244 : T241;
  assign T241 = T19 ? T243 : T242;
  assign T242 = io_in_acquire_bits_addr_block;
  assign T243 = io_in_acquire_bits_addr_block;
  assign T244 = io_in_acquire_bits_addr_block;
  assign T245 = io_in_acquire_bits_addr_block;
  assign T246 = R247;
  assign T248 = T88 ? io_in_acquire_bits_addr_block : R247;
  assign io_out_acquire_valid = T249;
  assign T249 = T251 | T250;
  assign T250 = T98 & ReorderQueue_io_enq_ready;
  assign T251 = R85 | T252;
  assign T252 = T254 & T253;
  assign T253 = T19 ^ 1'h1;
  assign T254 = io_in_acquire_valid & T255;
  assign T255 = T89 ^ 1'h1;
  assign io_in_grant_bits_data = T256;
  assign T256 = R105 ? T262 : T257;
  assign T257 = T77 ? T259 : T347;
  assign T347 = {64'h0, T258};
  assign T258 = io_out_grant_bits_data;
  assign T259 = T348;
  assign T348 = T260[7'h7f:1'h0];
  assign T260 = io_out_grant_bits_data << T261;
  assign T261 = {ReorderQueue_io_deq_data, 6'h0};
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = {R271, R265};
  assign T266 = T267 ? io_out_grant_bits_data : R265;
  assign T267 = T113 & T268;
  assign T268 = T269[1'h0];
  assign T269 = 1'h1 << T270;
  assign T270 = R110;
  assign T272 = T273 ? io_out_grant_bits_data : R271;
  assign T273 = T113 & T274;
  assign T274 = T269[1'h1];
  assign io_in_grant_bits_g_type = T275;
  assign T275 = R105 ? T279 : T276;
  assign T276 = T77 ? T278 : T277;
  assign T277 = io_out_grant_bits_g_type;
  assign T278 = 4'h4;
  assign T279 = 4'h5;
  assign io_in_grant_bits_is_builtin_type = T280;
  assign T280 = R105 ? T284 : T281;
  assign T281 = T77 ? T283 : T282;
  assign T282 = io_out_grant_bits_is_builtin_type;
  assign T283 = 1'h1;
  assign T284 = 1'h1;
  assign io_in_grant_bits_manager_xact_id = T285;
  assign T285 = R105 ? T289 : T286;
  assign T286 = T77 ? T288 : T287;
  assign T287 = io_out_grant_bits_manager_xact_id;
  assign T288 = io_out_grant_bits_manager_xact_id;
  assign T289 = R290;
  assign T291 = T108 ? io_out_grant_bits_manager_xact_id : R290;
  assign io_in_grant_bits_client_xact_id = T292;
  assign T292 = R105 ? T296 : T293;
  assign T293 = T77 ? T295 : T294;
  assign T294 = io_out_grant_bits_client_xact_id;
  assign T295 = io_out_grant_bits_client_xact_id;
  assign T296 = R297;
  assign T298 = T108 ? io_out_grant_bits_client_xact_id : R297;
  assign io_in_grant_bits_addr_beat = T349;
  assign T349 = T299[1'h1:1'h0];
  assign T299 = R105 ? T351 : T300;
  assign T300 = T77 ? T350 : T301;
  assign T301 = io_out_grant_bits_addr_beat;
  assign T350 = {1'h0, T302};
  assign T302 = T303;
  assign T303 = io_out_grant_bits_addr_beat >> 1'h1;
  assign T351 = {1'h0, T304};
  assign T304 = R305;
  assign T352 = reset ? 2'h0 : T306;
  assign T306 = T116 ? T307 : R305;
  assign T307 = R305 + 2'h1;
  assign io_in_grant_valid = T308;
  assign T308 = R105 | T309;
  assign T309 = io_out_grant_valid & T310;
  assign T310 = T101 ^ 1'h1;
  assign io_in_acquire_ready = T311;
  assign T311 = T317 & T312;
  assign T312 = T314 | T313;
  assign T313 = ReorderQueue_io_enq_ready & io_out_acquire_ready;
  assign T314 = T89 | T315;
  assign T315 = T316 & io_out_acquire_ready;
  assign T316 = T19 ^ 1'h1;
  assign T317 = R85 ^ 1'h1;
  ReorderQueue_0 ReorderQueue(.clk(clk), .reset(reset),
       .io_enq_ready( ReorderQueue_io_enq_ready ),
       .io_enq_valid( T83 ),
       .io_enq_bits_data( T79 ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T76 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( ReorderQueue_io_deq_data )
       //.io_deq_matches(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T21 <= 1'b1;
  if(!T22 && T21 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Put wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Get wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R85 <= 1'h0;
    end else if(T91) begin
      R85 <= 1'h0;
    end else if(T88) begin
      R85 <= 1'h1;
    end
    if(reset) begin
      R93 <= 1'h0;
    end else if(T96) begin
      R93 <= T95;
    end
    if(reset) begin
      R105 <= 1'h0;
    end else if(T116) begin
      R105 <= 1'h0;
    end else if(T108) begin
      R105 <= 1'h1;
    end
    if(reset) begin
      R110 <= 1'h0;
    end else if(T113) begin
      R110 <= T112;
    end
    if(T96) begin
      R135 <= T332;
    end else if(T88) begin
      R135 <= io_in_acquire_bits_data;
    end
    if(T96) begin
      R168 <= T343;
    end else if(T88) begin
      R168 <= T171;
    end
    if(T88) begin
      R225 <= io_in_acquire_bits_addr_beat;
    end
    if(T88) begin
      R236 <= io_in_acquire_bits_client_xact_id;
    end
    if(T88) begin
      R247 <= io_in_acquire_bits_addr_block;
    end
    if(T267) begin
      R265 <= io_out_grant_bits_data;
    end
    if(T273) begin
      R271 <= io_out_grant_bits_data;
    end
    if(T108) begin
      R290 <= io_out_grant_bits_manager_xact_id;
    end
    if(T108) begin
      R297 <= io_out_grant_bits_client_xact_id;
    end
    if(reset) begin
      R305 <= 2'h0;
    end else if(T116) begin
      R305 <= T307;
    end
  end
endmodule

module ReorderQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_data_addr_beat,
    input [2:0] io_enq_bits_data_byteOff,
    input  io_enq_bits_data_subblock,
    input [5:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [5:0] io_deq_tag,
    output[2:0] io_deq_data_addr_beat,
    output[2:0] io_deq_data_byteOff,
    output io_deq_data_subblock,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_8;
  wire T1;
  reg  roq_free_8;
  wire T250;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[15:0] T6;
  wire[3:0] T7;
  wire[3:0] roq_enq_addr;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  reg  roq_free_7;
  wire T251;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[15:0] T21;
  wire[3:0] T22;
  wire[3:0] roq_deq_addr;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire roq_matches_7;
  wire T30;
  wire T31;
  reg [5:0] roq_tags_7;
  wire[5:0] T32;
  wire T33;
  wire T34;
  wire[15:0] T35;
  wire[3:0] T36;
  wire roq_matches_6;
  wire T37;
  wire T38;
  reg [5:0] roq_tags_6;
  wire[5:0] T39;
  wire T40;
  wire T41;
  wire roq_matches_5;
  wire T42;
  wire T43;
  reg [5:0] roq_tags_5;
  wire[5:0] T44;
  wire T45;
  wire T46;
  wire roq_matches_4;
  wire T47;
  wire T48;
  reg [5:0] roq_tags_4;
  wire[5:0] T49;
  wire T50;
  wire T51;
  wire roq_matches_3;
  wire T52;
  wire T53;
  reg [5:0] roq_tags_3;
  wire[5:0] T54;
  wire T55;
  wire T56;
  wire roq_matches_2;
  wire T57;
  wire T58;
  reg [5:0] roq_tags_2;
  wire[5:0] T59;
  wire T60;
  wire T61;
  wire roq_matches_1;
  wire T62;
  wire T63;
  reg [5:0] roq_tags_1;
  wire[5:0] T64;
  wire T65;
  wire T66;
  wire roq_matches_0;
  wire T67;
  wire T68;
  reg [5:0] roq_tags_0;
  wire[5:0] T69;
  wire T70;
  wire T71;
  reg  roq_free_6;
  wire T252;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  roq_free_5;
  wire T253;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  reg  roq_free_4;
  wire T254;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  roq_free_3;
  wire T255;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  roq_free_2;
  wire T256;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  reg  roq_free_1;
  wire T257;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  roq_free_0;
  wire T258;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  reg [5:0] roq_tags_8;
  wire[5:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg  roq_data_0_subblock;
  wire T132;
  wire T133;
  wire T134;
  wire[15:0] T135;
  wire[3:0] T136;
  reg  roq_data_1_subblock;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  reg  roq_data_2_subblock;
  wire T143;
  wire T144;
  wire T145;
  reg  roq_data_3_subblock;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  roq_data_4_subblock;
  wire T153;
  wire T154;
  wire T155;
  reg  roq_data_5_subblock;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  reg  roq_data_6_subblock;
  wire T161;
  wire T162;
  wire T163;
  reg  roq_data_7_subblock;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  reg  roq_data_8_subblock;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire[2:0] T174;
  wire[2:0] T175;
  wire[2:0] T176;
  wire[2:0] T177;
  reg [2:0] roq_data_0_byteOff;
  wire[2:0] T178;
  wire T179;
  reg [2:0] roq_data_1_byteOff;
  wire[2:0] T180;
  wire T181;
  wire T182;
  wire[2:0] T183;
  reg [2:0] roq_data_2_byteOff;
  wire[2:0] T184;
  wire T185;
  reg [2:0] roq_data_3_byteOff;
  wire[2:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire[2:0] T190;
  wire[2:0] T191;
  reg [2:0] roq_data_4_byteOff;
  wire[2:0] T192;
  wire T193;
  reg [2:0] roq_data_5_byteOff;
  wire[2:0] T194;
  wire T195;
  wire T196;
  wire[2:0] T197;
  reg [2:0] roq_data_6_byteOff;
  wire[2:0] T198;
  wire T199;
  reg [2:0] roq_data_7_byteOff;
  wire[2:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  reg [2:0] roq_data_8_byteOff;
  wire[2:0] T205;
  wire T206;
  wire T207;
  wire[2:0] T208;
  wire[2:0] T209;
  wire[2:0] T210;
  wire[2:0] T211;
  reg [2:0] roq_data_0_addr_beat;
  wire[2:0] T212;
  wire T213;
  reg [2:0] roq_data_1_addr_beat;
  wire[2:0] T214;
  wire T215;
  wire T216;
  wire[2:0] T217;
  reg [2:0] roq_data_2_addr_beat;
  wire[2:0] T218;
  wire T219;
  reg [2:0] roq_data_3_addr_beat;
  wire[2:0] T220;
  wire T221;
  wire T222;
  wire T223;
  wire[2:0] T224;
  wire[2:0] T225;
  reg [2:0] roq_data_4_addr_beat;
  wire[2:0] T226;
  wire T227;
  reg [2:0] roq_data_5_addr_beat;
  wire[2:0] T228;
  wire T229;
  wire T230;
  wire[2:0] T231;
  reg [2:0] roq_data_6_addr_beat;
  wire[2:0] T232;
  wire T233;
  reg [2:0] roq_data_7_addr_beat;
  wire[2:0] T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  reg [2:0] roq_data_8_addr_beat;
  wire[2:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_8 = {1{$random}};
    roq_free_7 = {1{$random}};
    roq_tags_7 = {1{$random}};
    roq_tags_6 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_6 = {1{$random}};
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_8 = {1{$random}};
    roq_data_0_subblock = {1{$random}};
    roq_data_1_subblock = {1{$random}};
    roq_data_2_subblock = {1{$random}};
    roq_data_3_subblock = {1{$random}};
    roq_data_4_subblock = {1{$random}};
    roq_data_5_subblock = {1{$random}};
    roq_data_6_subblock = {1{$random}};
    roq_data_7_subblock = {1{$random}};
    roq_data_8_subblock = {1{$random}};
    roq_data_0_byteOff = {1{$random}};
    roq_data_1_byteOff = {1{$random}};
    roq_data_2_byteOff = {1{$random}};
    roq_data_3_byteOff = {1{$random}};
    roq_data_4_byteOff = {1{$random}};
    roq_data_5_byteOff = {1{$random}};
    roq_data_6_byteOff = {1{$random}};
    roq_data_7_byteOff = {1{$random}};
    roq_data_8_byteOff = {1{$random}};
    roq_data_0_addr_beat = {1{$random}};
    roq_data_1_addr_beat = {1{$random}};
    roq_data_2_addr_beat = {1{$random}};
    roq_data_3_addr_beat = {1{$random}};
    roq_data_4_addr_beat = {1{$random}};
    roq_data_5_addr_beat = {1{$random}};
    roq_data_6_addr_beat = {1{$random}};
    roq_data_7_addr_beat = {1{$random}};
    roq_data_8_addr_beat = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T121 | roq_matches_8;
  assign roq_matches_8 = T117 & T1;
  assign T1 = roq_free_8 ^ 1'h1;
  assign T250 = reset ? 1'h1 : T2;
  assign T2 = T115 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_8;
  assign T4 = T114 & T5;
  assign T5 = T6[4'h8];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 4'h0 : T8;
  assign T8 = roq_free_1 ? 4'h1 : T9;
  assign T9 = roq_free_2 ? 4'h2 : T10;
  assign T10 = roq_free_3 ? 4'h3 : T11;
  assign T11 = roq_free_4 ? 4'h4 : T12;
  assign T12 = roq_free_5 ? 4'h5 : T13;
  assign T13 = roq_free_6 ? 4'h6 : T14;
  assign T14 = roq_free_7 ? 4'h7 : 4'h8;
  assign T251 = reset ? 1'h1 : T15;
  assign T15 = T19 ? 1'h1 : T16;
  assign T16 = T17 ? 1'h0 : roq_free_7;
  assign T17 = T114 & T18;
  assign T18 = T6[3'h7];
  assign T19 = io_deq_valid & T20;
  assign T20 = T21[3'h7];
  assign T21 = 1'h1 << T22;
  assign T22 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 4'h0 : T23;
  assign T23 = roq_matches_1 ? 4'h1 : T24;
  assign T24 = roq_matches_2 ? 4'h2 : T25;
  assign T25 = roq_matches_3 ? 4'h3 : T26;
  assign T26 = roq_matches_4 ? 4'h4 : T27;
  assign T27 = roq_matches_5 ? 4'h5 : T28;
  assign T28 = roq_matches_6 ? 4'h6 : T29;
  assign T29 = roq_matches_7 ? 4'h7 : 4'h8;
  assign roq_matches_7 = T31 & T30;
  assign T30 = roq_free_7 ^ 1'h1;
  assign T31 = roq_tags_7 == io_deq_tag;
  assign T32 = T33 ? io_enq_bits_tag : roq_tags_7;
  assign T33 = T114 & T34;
  assign T34 = T35[3'h7];
  assign T35 = 1'h1 << T36;
  assign T36 = roq_enq_addr;
  assign roq_matches_6 = T38 & T37;
  assign T37 = roq_free_6 ^ 1'h1;
  assign T38 = roq_tags_6 == io_deq_tag;
  assign T39 = T40 ? io_enq_bits_tag : roq_tags_6;
  assign T40 = T114 & T41;
  assign T41 = T35[3'h6];
  assign roq_matches_5 = T43 & T42;
  assign T42 = roq_free_5 ^ 1'h1;
  assign T43 = roq_tags_5 == io_deq_tag;
  assign T44 = T45 ? io_enq_bits_tag : roq_tags_5;
  assign T45 = T114 & T46;
  assign T46 = T35[3'h5];
  assign roq_matches_4 = T48 & T47;
  assign T47 = roq_free_4 ^ 1'h1;
  assign T48 = roq_tags_4 == io_deq_tag;
  assign T49 = T50 ? io_enq_bits_tag : roq_tags_4;
  assign T50 = T114 & T51;
  assign T51 = T35[3'h4];
  assign roq_matches_3 = T53 & T52;
  assign T52 = roq_free_3 ^ 1'h1;
  assign T53 = roq_tags_3 == io_deq_tag;
  assign T54 = T55 ? io_enq_bits_tag : roq_tags_3;
  assign T55 = T114 & T56;
  assign T56 = T35[2'h3];
  assign roq_matches_2 = T58 & T57;
  assign T57 = roq_free_2 ^ 1'h1;
  assign T58 = roq_tags_2 == io_deq_tag;
  assign T59 = T60 ? io_enq_bits_tag : roq_tags_2;
  assign T60 = T114 & T61;
  assign T61 = T35[2'h2];
  assign roq_matches_1 = T63 & T62;
  assign T62 = roq_free_1 ^ 1'h1;
  assign T63 = roq_tags_1 == io_deq_tag;
  assign T64 = T65 ? io_enq_bits_tag : roq_tags_1;
  assign T65 = T114 & T66;
  assign T66 = T35[1'h1];
  assign roq_matches_0 = T68 & T67;
  assign T67 = roq_free_0 ^ 1'h1;
  assign T68 = roq_tags_0 == io_deq_tag;
  assign T69 = T70 ? io_enq_bits_tag : roq_tags_0;
  assign T70 = T114 & T71;
  assign T71 = T35[1'h0];
  assign T252 = reset ? 1'h1 : T72;
  assign T72 = T76 ? 1'h1 : T73;
  assign T73 = T74 ? 1'h0 : roq_free_6;
  assign T74 = T114 & T75;
  assign T75 = T6[3'h6];
  assign T76 = io_deq_valid & T77;
  assign T77 = T21[3'h6];
  assign T253 = reset ? 1'h1 : T78;
  assign T78 = T82 ? 1'h1 : T79;
  assign T79 = T80 ? 1'h0 : roq_free_5;
  assign T80 = T114 & T81;
  assign T81 = T6[3'h5];
  assign T82 = io_deq_valid & T83;
  assign T83 = T21[3'h5];
  assign T254 = reset ? 1'h1 : T84;
  assign T84 = T88 ? 1'h1 : T85;
  assign T85 = T86 ? 1'h0 : roq_free_4;
  assign T86 = T114 & T87;
  assign T87 = T6[3'h4];
  assign T88 = io_deq_valid & T89;
  assign T89 = T21[3'h4];
  assign T255 = reset ? 1'h1 : T90;
  assign T90 = T94 ? 1'h1 : T91;
  assign T91 = T92 ? 1'h0 : roq_free_3;
  assign T92 = T114 & T93;
  assign T93 = T6[2'h3];
  assign T94 = io_deq_valid & T95;
  assign T95 = T21[2'h3];
  assign T256 = reset ? 1'h1 : T96;
  assign T96 = T100 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : roq_free_2;
  assign T98 = T114 & T99;
  assign T99 = T6[2'h2];
  assign T100 = io_deq_valid & T101;
  assign T101 = T21[2'h2];
  assign T257 = reset ? 1'h1 : T102;
  assign T102 = T106 ? 1'h1 : T103;
  assign T103 = T104 ? 1'h0 : roq_free_1;
  assign T104 = T114 & T105;
  assign T105 = T6[1'h1];
  assign T106 = io_deq_valid & T107;
  assign T107 = T21[1'h1];
  assign T258 = reset ? 1'h1 : T108;
  assign T108 = T112 ? 1'h1 : T109;
  assign T109 = T110 ? 1'h0 : roq_free_0;
  assign T110 = T114 & T111;
  assign T111 = T6[1'h0];
  assign T112 = io_deq_valid & T113;
  assign T113 = T21[1'h0];
  assign T114 = io_enq_valid & io_enq_ready;
  assign T115 = io_deq_valid & T116;
  assign T116 = T21[4'h8];
  assign T117 = roq_tags_8 == io_deq_tag;
  assign T118 = T119 ? io_enq_bits_tag : roq_tags_8;
  assign T119 = T114 & T120;
  assign T120 = T35[4'h8];
  assign T121 = T122 | roq_matches_7;
  assign T122 = T123 | roq_matches_6;
  assign T123 = T124 | roq_matches_5;
  assign T124 = T125 | roq_matches_4;
  assign T125 = T126 | roq_matches_3;
  assign T126 = T127 | roq_matches_2;
  assign T127 = roq_matches_0 | roq_matches_1;
  assign io_deq_data_subblock = T128;
  assign T128 = T173 ? roq_data_8_subblock : T129;
  assign T129 = T169 ? T151 : T130;
  assign T130 = T150 ? T142 : T131;
  assign T131 = T140 ? roq_data_1_subblock : roq_data_0_subblock;
  assign T132 = T133 ? io_enq_bits_data_subblock : roq_data_0_subblock;
  assign T133 = T114 & T134;
  assign T134 = T135[1'h0];
  assign T135 = 1'h1 << T136;
  assign T136 = roq_enq_addr;
  assign T137 = T138 ? io_enq_bits_data_subblock : roq_data_1_subblock;
  assign T138 = T114 & T139;
  assign T139 = T135[1'h1];
  assign T140 = T141[1'h0];
  assign T141 = roq_deq_addr;
  assign T142 = T149 ? roq_data_3_subblock : roq_data_2_subblock;
  assign T143 = T144 ? io_enq_bits_data_subblock : roq_data_2_subblock;
  assign T144 = T114 & T145;
  assign T145 = T135[2'h2];
  assign T146 = T147 ? io_enq_bits_data_subblock : roq_data_3_subblock;
  assign T147 = T114 & T148;
  assign T148 = T135[2'h3];
  assign T149 = T141[1'h0];
  assign T150 = T141[1'h1];
  assign T151 = T168 ? T160 : T152;
  assign T152 = T159 ? roq_data_5_subblock : roq_data_4_subblock;
  assign T153 = T154 ? io_enq_bits_data_subblock : roq_data_4_subblock;
  assign T154 = T114 & T155;
  assign T155 = T135[3'h4];
  assign T156 = T157 ? io_enq_bits_data_subblock : roq_data_5_subblock;
  assign T157 = T114 & T158;
  assign T158 = T135[3'h5];
  assign T159 = T141[1'h0];
  assign T160 = T167 ? roq_data_7_subblock : roq_data_6_subblock;
  assign T161 = T162 ? io_enq_bits_data_subblock : roq_data_6_subblock;
  assign T162 = T114 & T163;
  assign T163 = T135[3'h6];
  assign T164 = T165 ? io_enq_bits_data_subblock : roq_data_7_subblock;
  assign T165 = T114 & T166;
  assign T166 = T135[3'h7];
  assign T167 = T141[1'h0];
  assign T168 = T141[1'h1];
  assign T169 = T141[2'h2];
  assign T170 = T171 ? io_enq_bits_data_subblock : roq_data_8_subblock;
  assign T171 = T114 & T172;
  assign T172 = T135[4'h8];
  assign T173 = T141[2'h3];
  assign io_deq_data_byteOff = T174;
  assign T174 = T207 ? roq_data_8_byteOff : T175;
  assign T175 = T204 ? T190 : T176;
  assign T176 = T189 ? T183 : T177;
  assign T177 = T182 ? roq_data_1_byteOff : roq_data_0_byteOff;
  assign T178 = T179 ? io_enq_bits_data_byteOff : roq_data_0_byteOff;
  assign T179 = T114 & T134;
  assign T180 = T181 ? io_enq_bits_data_byteOff : roq_data_1_byteOff;
  assign T181 = T114 & T139;
  assign T182 = T141[1'h0];
  assign T183 = T188 ? roq_data_3_byteOff : roq_data_2_byteOff;
  assign T184 = T185 ? io_enq_bits_data_byteOff : roq_data_2_byteOff;
  assign T185 = T114 & T145;
  assign T186 = T187 ? io_enq_bits_data_byteOff : roq_data_3_byteOff;
  assign T187 = T114 & T148;
  assign T188 = T141[1'h0];
  assign T189 = T141[1'h1];
  assign T190 = T203 ? T197 : T191;
  assign T191 = T196 ? roq_data_5_byteOff : roq_data_4_byteOff;
  assign T192 = T193 ? io_enq_bits_data_byteOff : roq_data_4_byteOff;
  assign T193 = T114 & T155;
  assign T194 = T195 ? io_enq_bits_data_byteOff : roq_data_5_byteOff;
  assign T195 = T114 & T158;
  assign T196 = T141[1'h0];
  assign T197 = T202 ? roq_data_7_byteOff : roq_data_6_byteOff;
  assign T198 = T199 ? io_enq_bits_data_byteOff : roq_data_6_byteOff;
  assign T199 = T114 & T163;
  assign T200 = T201 ? io_enq_bits_data_byteOff : roq_data_7_byteOff;
  assign T201 = T114 & T166;
  assign T202 = T141[1'h0];
  assign T203 = T141[1'h1];
  assign T204 = T141[2'h2];
  assign T205 = T206 ? io_enq_bits_data_byteOff : roq_data_8_byteOff;
  assign T206 = T114 & T172;
  assign T207 = T141[2'h3];
  assign io_deq_data_addr_beat = T208;
  assign T208 = T241 ? roq_data_8_addr_beat : T209;
  assign T209 = T238 ? T224 : T210;
  assign T210 = T223 ? T217 : T211;
  assign T211 = T216 ? roq_data_1_addr_beat : roq_data_0_addr_beat;
  assign T212 = T213 ? io_enq_bits_data_addr_beat : roq_data_0_addr_beat;
  assign T213 = T114 & T134;
  assign T214 = T215 ? io_enq_bits_data_addr_beat : roq_data_1_addr_beat;
  assign T215 = T114 & T139;
  assign T216 = T141[1'h0];
  assign T217 = T222 ? roq_data_3_addr_beat : roq_data_2_addr_beat;
  assign T218 = T219 ? io_enq_bits_data_addr_beat : roq_data_2_addr_beat;
  assign T219 = T114 & T145;
  assign T220 = T221 ? io_enq_bits_data_addr_beat : roq_data_3_addr_beat;
  assign T221 = T114 & T148;
  assign T222 = T141[1'h0];
  assign T223 = T141[1'h1];
  assign T224 = T237 ? T231 : T225;
  assign T225 = T230 ? roq_data_5_addr_beat : roq_data_4_addr_beat;
  assign T226 = T227 ? io_enq_bits_data_addr_beat : roq_data_4_addr_beat;
  assign T227 = T114 & T155;
  assign T228 = T229 ? io_enq_bits_data_addr_beat : roq_data_5_addr_beat;
  assign T229 = T114 & T158;
  assign T230 = T141[1'h0];
  assign T231 = T236 ? roq_data_7_addr_beat : roq_data_6_addr_beat;
  assign T232 = T233 ? io_enq_bits_data_addr_beat : roq_data_6_addr_beat;
  assign T233 = T114 & T163;
  assign T234 = T235 ? io_enq_bits_data_addr_beat : roq_data_7_addr_beat;
  assign T235 = T114 & T166;
  assign T236 = T141[1'h0];
  assign T237 = T141[1'h1];
  assign T238 = T141[2'h2];
  assign T239 = T240 ? io_enq_bits_data_addr_beat : roq_data_8_addr_beat;
  assign T240 = T114 & T172;
  assign T241 = T141[2'h3];
  assign io_enq_ready = T242;
  assign T242 = T243 | roq_free_8;
  assign T243 = T244 | roq_free_7;
  assign T244 = T245 | roq_free_6;
  assign T245 = T246 | roq_free_5;
  assign T246 = T247 | roq_free_4;
  assign T247 = T248 | roq_free_3;
  assign T248 = T249 | roq_free_2;
  assign T249 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_8 <= 1'h1;
    end else if(T115) begin
      roq_free_8 <= 1'h1;
    end else if(T4) begin
      roq_free_8 <= 1'h0;
    end
    if(reset) begin
      roq_free_7 <= 1'h1;
    end else if(T19) begin
      roq_free_7 <= 1'h1;
    end else if(T17) begin
      roq_free_7 <= 1'h0;
    end
    if(T33) begin
      roq_tags_7 <= io_enq_bits_tag;
    end
    if(T40) begin
      roq_tags_6 <= io_enq_bits_tag;
    end
    if(T45) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T50) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T55) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T60) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T65) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T70) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_6 <= 1'h1;
    end else if(T76) begin
      roq_free_6 <= 1'h1;
    end else if(T74) begin
      roq_free_6 <= 1'h0;
    end
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T82) begin
      roq_free_5 <= 1'h1;
    end else if(T80) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T88) begin
      roq_free_4 <= 1'h1;
    end else if(T86) begin
      roq_free_4 <= 1'h0;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T94) begin
      roq_free_3 <= 1'h1;
    end else if(T92) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T100) begin
      roq_free_2 <= 1'h1;
    end else if(T98) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T106) begin
      roq_free_1 <= 1'h1;
    end else if(T104) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T112) begin
      roq_free_0 <= 1'h1;
    end else if(T110) begin
      roq_free_0 <= 1'h0;
    end
    if(T119) begin
      roq_tags_8 <= io_enq_bits_tag;
    end
    if(T133) begin
      roq_data_0_subblock <= io_enq_bits_data_subblock;
    end
    if(T138) begin
      roq_data_1_subblock <= io_enq_bits_data_subblock;
    end
    if(T144) begin
      roq_data_2_subblock <= io_enq_bits_data_subblock;
    end
    if(T147) begin
      roq_data_3_subblock <= io_enq_bits_data_subblock;
    end
    if(T154) begin
      roq_data_4_subblock <= io_enq_bits_data_subblock;
    end
    if(T157) begin
      roq_data_5_subblock <= io_enq_bits_data_subblock;
    end
    if(T162) begin
      roq_data_6_subblock <= io_enq_bits_data_subblock;
    end
    if(T165) begin
      roq_data_7_subblock <= io_enq_bits_data_subblock;
    end
    if(T171) begin
      roq_data_8_subblock <= io_enq_bits_data_subblock;
    end
    if(T179) begin
      roq_data_0_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T181) begin
      roq_data_1_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T185) begin
      roq_data_2_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T187) begin
      roq_data_3_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T193) begin
      roq_data_4_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T195) begin
      roq_data_5_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T199) begin
      roq_data_6_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T201) begin
      roq_data_7_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T206) begin
      roq_data_8_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T213) begin
      roq_data_0_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T215) begin
      roq_data_1_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T219) begin
      roq_data_2_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T221) begin
      roq_data_3_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T227) begin
      roq_data_4_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T229) begin
      roq_data_5_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T233) begin
      roq_data_6_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T235) begin
      roq_data_7_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T240) begin
      roq_data_8_addr_beat <= io_enq_bits_data_addr_beat;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_addr_beat,
    input [3:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_addr_beat,
    input [3:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_addr_beat,
    output[3:0] io_out_bits_client_xact_id,
    output io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[63:0] io_out_bits_data,
    output io_out_bits_client_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[3:0] T3;
  wire T4;
  wire T5;
  wire[3:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_client_id = T0;
  assign T0 = T1 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_g_type = T3;
  assign T3 = T1 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign io_out_bits_is_builtin_type = T4;
  assign T4 = T1 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module NastiIOTileLinkIOConverter(input clk, input reset,
    output io_tl_acquire_ready,
    input  io_tl_acquire_valid,
    input [25:0] io_tl_acquire_bits_addr_block,
    input [3:0] io_tl_acquire_bits_client_xact_id,
    input [2:0] io_tl_acquire_bits_addr_beat,
    input  io_tl_acquire_bits_is_builtin_type,
    input [2:0] io_tl_acquire_bits_a_type,
    input [11:0] io_tl_acquire_bits_union,
    input [63:0] io_tl_acquire_bits_data,
    input  io_tl_grant_ready,
    output io_tl_grant_valid,
    output[2:0] io_tl_grant_bits_addr_beat,
    output[3:0] io_tl_grant_bits_client_xact_id,
    output io_tl_grant_bits_manager_xact_id,
    output io_tl_grant_bits_is_builtin_type,
    output[3:0] io_tl_grant_bits_g_type,
    output[63:0] io_tl_grant_bits_data,
    input  io_nasti_aw_ready,
    output io_nasti_aw_valid,
    output[31:0] io_nasti_aw_bits_addr,
    output[7:0] io_nasti_aw_bits_len,
    output[2:0] io_nasti_aw_bits_size,
    output[1:0] io_nasti_aw_bits_burst,
    output io_nasti_aw_bits_lock,
    output[3:0] io_nasti_aw_bits_cache,
    output[2:0] io_nasti_aw_bits_prot,
    output[3:0] io_nasti_aw_bits_qos,
    output[3:0] io_nasti_aw_bits_region,
    output[5:0] io_nasti_aw_bits_id,
    output io_nasti_aw_bits_user,
    input  io_nasti_w_ready,
    output io_nasti_w_valid,
    output[63:0] io_nasti_w_bits_data,
    output io_nasti_w_bits_last,
    output[7:0] io_nasti_w_bits_strb,
    output io_nasti_w_bits_user,
    output io_nasti_b_ready,
    input  io_nasti_b_valid,
    input [1:0] io_nasti_b_bits_resp,
    input [5:0] io_nasti_b_bits_id,
    input  io_nasti_b_bits_user,
    input  io_nasti_ar_ready,
    output io_nasti_ar_valid,
    output[31:0] io_nasti_ar_bits_addr,
    output[7:0] io_nasti_ar_bits_len,
    output[2:0] io_nasti_ar_bits_size,
    output[1:0] io_nasti_ar_bits_burst,
    output io_nasti_ar_bits_lock,
    output[3:0] io_nasti_ar_bits_cache,
    output[2:0] io_nasti_ar_bits_prot,
    output[3:0] io_nasti_ar_bits_qos,
    output[3:0] io_nasti_ar_bits_region,
    output[5:0] io_nasti_ar_bits_id,
    output io_nasti_ar_bits_user,
    output io_nasti_r_ready,
    input  io_nasti_r_valid,
    input [1:0] io_nasti_r_bits_resp,
    input [63:0] io_nasti_r_bits_data,
    input  io_nasti_r_bits_last,
    input [5:0] io_nasti_r_bits_id,
    input  io_nasti_r_bits_user
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg  T10;
  wire T11;
  wire T12;
  wire T13;
  wire[63:0] T14;
  wire[63:0] T146;
  wire[126:0] r_aligned_data;
  wire[126:0] T147;
  wire[126:0] T15;
  wire[5:0] T16;
  wire[3:0] T17;
  wire[3:0] T148;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T149;
  wire[2:0] T22;
  wire[2:0] T23;
  reg [2:0] tl_cnt_in;
  wire[2:0] T150;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[63:0] T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire[3:0] T35;
  wire[3:0] T151;
  wire[2:0] T36;
  wire T37;
  wire T38;
  wire nasti_wrap_out;
  wire T39;
  reg [2:0] nasti_cnt_out;
  wire[2:0] T152;
  wire[2:0] T40;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire is_subblock;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire get_valid;
  wire T53;
  wire has_data;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire[5:0] T60;
  wire[5:0] T153;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[2:0] T63;
  wire[3:0] T64;
  wire T65;
  wire[1:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire[7:0] T154;
  wire[2:0] T87;
  wire[31:0] T88;
  wire[31:0] T89;
  wire[5:0] T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire[7:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[7:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire tl_wrap_out;
  wire T110;
  reg [2:0] tl_cnt_out;
  wire[2:0] T155;
  wire[2:0] T111;
  wire[2:0] T112;
  wire T113;
  wire is_multibeat;
  wire T114;
  wire T115;
  wire[63:0] T116;
  wire T117;
  wire aw_ready;
  reg  w_inflight;
  wire T156;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire put_valid;
  wire T125;
  wire[5:0] T126;
  wire[5:0] T157;
  wire[3:0] T127;
  wire[3:0] T128;
  wire[2:0] T129;
  wire[3:0] T130;
  wire T131;
  wire[1:0] T132;
  wire[2:0] T133;
  wire[7:0] T134;
  wire[7:0] T158;
  wire[2:0] T135;
  wire[31:0] T136;
  wire[31:0] T137;
  wire[5:0] T138;
  wire[2:0] T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire roq_io_enq_ready;
  wire[2:0] roq_io_deq_data_addr_beat;
  wire[2:0] roq_io_deq_data_byteOff;
  wire roq_io_deq_data_subblock;
  wire roq_io_deq_matches;
  wire gnt_arb_io_in_1_ready;
  wire gnt_arb_io_in_0_ready;
  wire gnt_arb_io_out_valid;
  wire[2:0] gnt_arb_io_out_bits_addr_beat;
  wire[3:0] gnt_arb_io_out_bits_client_xact_id;
  wire gnt_arb_io_out_bits_manager_xact_id;
  wire gnt_arb_io_out_bits_is_builtin_type;
  wire[3:0] gnt_arb_io_out_bits_g_type;
  wire[63:0] gnt_arb_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T5 = 1'b0;
    T10 = 1'b0;
    tl_cnt_in = {1{$random}};
    nasti_cnt_out = {1{$random}};
    tl_cnt_out = {1{$random}};
    w_inflight = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = io_nasti_b_bits_resp == 2'h0;
  assign T4 = io_nasti_b_valid ^ 1'h1;
  assign T6 = T7 | reset;
  assign T7 = T9 | T8;
  assign T8 = io_nasti_r_bits_resp == 2'h0;
  assign T9 = io_nasti_r_valid ^ 1'h1;
  assign T11 = T12 | reset;
  assign T12 = T13 | roq_io_deq_matches;
  assign T13 = io_nasti_r_valid ^ 1'h1;
  assign T14 = T146;
  assign T146 = r_aligned_data[6'h3f:1'h0];
  assign r_aligned_data = roq_io_deq_data_subblock ? T15 : T147;
  assign T147 = {63'h0, io_nasti_r_bits_data};
  assign T15 = io_nasti_r_bits_data << T16;
  assign T16 = {roq_io_deq_data_byteOff, 3'h0};
  assign T17 = T148;
  assign T148 = {1'h0, T18};
  assign T18 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T19 = 1'h1;
  assign T20 = 1'h0;
  assign T21 = T149;
  assign T149 = io_nasti_r_bits_id[2'h3:1'h0];
  assign T22 = T23;
  assign T23 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T150 = reset ? 3'h0 : T24;
  assign T24 = T26 ? T25 : tl_cnt_in;
  assign T25 = tl_cnt_in + 3'h1;
  assign T26 = T30 & T27;
  assign T27 = io_tl_grant_bits_is_builtin_type ? T29 : T28;
  assign T28 = 4'h0 == io_tl_grant_bits_g_type;
  assign T29 = 4'h5 == io_tl_grant_bits_g_type;
  assign T30 = io_tl_grant_ready & io_tl_grant_valid;
  assign T31 = 64'h0;
  assign T32 = 4'h3;
  assign T33 = 1'h1;
  assign T34 = 1'h0;
  assign T35 = T151;
  assign T151 = io_nasti_b_bits_id[2'h3:1'h0];
  assign T36 = 3'h0;
  assign T37 = T45 & T38;
  assign T38 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign nasti_wrap_out = T42 & T39;
  assign T39 = nasti_cnt_out == 3'h7;
  assign T152 = reset ? 3'h0 : T40;
  assign T40 = T42 ? T41 : nasti_cnt_out;
  assign T41 = nasti_cnt_out + 3'h1;
  assign T42 = T44 & T43;
  assign T43 = roq_io_deq_data_subblock ^ 1'h1;
  assign T44 = io_nasti_r_ready & io_nasti_r_valid;
  assign T45 = io_nasti_r_ready & io_nasti_r_valid;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T46;
  assign T46 = T48 | T47;
  assign T47 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T48 = T50 | T49;
  assign T49 = 3'h0 == io_tl_acquire_bits_a_type;
  assign T50 = 3'h2 == io_tl_acquire_bits_a_type;
  assign T51 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign T52 = get_valid & io_nasti_ar_ready;
  assign get_valid = io_tl_acquire_valid & T53;
  assign T53 = has_data ^ 1'h1;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T54;
  assign T54 = T56 | T55;
  assign T55 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T56 = T58 | T57;
  assign T57 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T58 = 3'h2 == io_tl_acquire_bits_a_type;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign io_nasti_ar_bits_user = T59;
  assign T59 = 1'h0;
  assign io_nasti_ar_bits_id = T60;
  assign T60 = T153;
  assign T153 = {2'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_ar_bits_region = T61;
  assign T61 = 4'h0;
  assign io_nasti_ar_bits_qos = T62;
  assign T62 = 4'h0;
  assign io_nasti_ar_bits_prot = T63;
  assign T63 = 3'h0;
  assign io_nasti_ar_bits_cache = T64;
  assign T64 = 4'h0;
  assign io_nasti_ar_bits_lock = T65;
  assign T65 = 1'h0;
  assign io_nasti_ar_bits_burst = T66;
  assign T66 = 2'h1;
  assign io_nasti_ar_bits_size = T67;
  assign T67 = T68;
  assign T68 = is_subblock ? T69 : 3'h3;
  assign T69 = T85 ? 3'h0 : T70;
  assign T70 = T84 ? 3'h0 : T71;
  assign T71 = T83 ? 3'h1 : T72;
  assign T72 = T82 ? 3'h1 : T73;
  assign T73 = T81 ? 3'h2 : T74;
  assign T74 = T80 ? 3'h2 : T75;
  assign T75 = T79 ? 3'h3 : T76;
  assign T76 = T77 ? 3'h3 : 3'h7;
  assign T77 = T78 == 3'h7;
  assign T78 = io_tl_acquire_bits_union[4'h8:3'h6];
  assign T79 = T78 == 3'h3;
  assign T80 = T78 == 3'h6;
  assign T81 = T78 == 3'h2;
  assign T82 = T78 == 3'h5;
  assign T83 = T78 == 3'h1;
  assign T84 = T78 == 3'h4;
  assign T85 = T78 == 3'h0;
  assign io_nasti_ar_bits_len = T86;
  assign T86 = T154;
  assign T154 = {5'h0, T87};
  assign T87 = is_subblock ? 3'h0 : 3'h7;
  assign io_nasti_ar_bits_addr = T88;
  assign T88 = T89;
  assign T89 = {io_tl_acquire_bits_addr_block, T90};
  assign T90 = {io_tl_acquire_bits_addr_beat, T91};
  assign T91 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_ar_valid = T92;
  assign T92 = get_valid & roq_io_enq_ready;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_w_bits_user = T93;
  assign T93 = 1'h0;
  assign io_nasti_w_bits_strb = T94;
  assign T94 = T95;
  assign T95 = T104 ? T103 : T96;
  assign T96 = T98 ? T97 : 8'h0;
  assign T97 = io_tl_acquire_bits_union[4'h8:1'h1];
  assign T98 = T101 | T99;
  assign T99 = io_tl_acquire_bits_is_builtin_type & T100;
  assign T100 = io_tl_acquire_bits_a_type == 3'h2;
  assign T101 = io_tl_acquire_bits_is_builtin_type & T102;
  assign T102 = io_tl_acquire_bits_a_type == 3'h3;
  assign T103 = 8'hff;
  assign T104 = io_tl_acquire_bits_is_builtin_type & T105;
  assign T105 = io_tl_acquire_bits_a_type == 3'h4;
  assign io_nasti_w_bits_last = T106;
  assign T106 = T107;
  assign T107 = tl_wrap_out | T108;
  assign T108 = T109 & is_subblock;
  assign T109 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign tl_wrap_out = T113 & T110;
  assign T110 = tl_cnt_out == 3'h7;
  assign T155 = reset ? 3'h0 : T111;
  assign T111 = T113 ? T112 : tl_cnt_out;
  assign T112 = tl_cnt_out + 3'h1;
  assign T113 = T115 & is_multibeat;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T114;
  assign T114 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T115 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign io_nasti_w_bits_data = T116;
  assign T116 = io_tl_acquire_bits_data;
  assign io_nasti_w_valid = T117;
  assign T117 = put_valid & aw_ready;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T156 = reset ? 1'h0 : T118;
  assign T118 = T124 ? 1'h0 : T119;
  assign T119 = T120 ? 1'h1 : w_inflight;
  assign T120 = T121 & is_multibeat;
  assign T121 = T123 & T122;
  assign T122 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T123 = w_inflight ^ 1'h1;
  assign T124 = w_inflight & tl_wrap_out;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign io_nasti_aw_bits_user = T125;
  assign T125 = 1'h0;
  assign io_nasti_aw_bits_id = T126;
  assign T126 = T157;
  assign T157 = {2'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_aw_bits_region = T127;
  assign T127 = 4'h0;
  assign io_nasti_aw_bits_qos = T128;
  assign T128 = 4'h0;
  assign io_nasti_aw_bits_prot = T129;
  assign T129 = 3'h0;
  assign io_nasti_aw_bits_cache = T130;
  assign T130 = 4'h0;
  assign io_nasti_aw_bits_lock = T131;
  assign T131 = 1'h0;
  assign io_nasti_aw_bits_burst = T132;
  assign T132 = 2'h1;
  assign io_nasti_aw_bits_size = T133;
  assign T133 = 3'h3;
  assign io_nasti_aw_bits_len = T134;
  assign T134 = T158;
  assign T158 = {5'h0, T135};
  assign T135 = is_multibeat ? 3'h7 : 3'h0;
  assign io_nasti_aw_bits_addr = T136;
  assign T136 = T137;
  assign T137 = {io_tl_acquire_bits_addr_block, T138};
  assign T138 = {io_tl_acquire_bits_addr_beat, T139};
  assign T139 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_aw_valid = T140;
  assign T140 = T142 & T141;
  assign T141 = w_inflight ^ 1'h1;
  assign T142 = put_valid & io_nasti_w_ready;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_acquire_ready = T143;
  assign T143 = has_data ? T145 : T144;
  assign T144 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T145 = aw_ready & io_nasti_w_ready;
  ReorderQueue_1 roq(.clk(clk), .reset(reset),
       .io_enq_ready( roq_io_enq_ready ),
       .io_enq_valid( T52 ),
       .io_enq_bits_data_addr_beat( io_tl_acquire_bits_addr_beat ),
       .io_enq_bits_data_byteOff( T51 ),
       .io_enq_bits_data_subblock( is_subblock ),
       .io_enq_bits_tag( io_nasti_ar_bits_id ),
       .io_deq_valid( T37 ),
       .io_deq_tag( io_nasti_r_bits_id ),
       .io_deq_data_addr_beat( roq_io_deq_data_addr_beat ),
       .io_deq_data_byteOff( roq_io_deq_data_byteOff ),
       .io_deq_data_subblock( roq_io_deq_data_subblock ),
       .io_deq_matches( roq_io_deq_matches )
  );
  Arbiter_6 gnt_arb(
       .io_in_1_ready( gnt_arb_io_in_1_ready ),
       .io_in_1_valid( io_nasti_b_valid ),
       .io_in_1_bits_addr_beat( T36 ),
       .io_in_1_bits_client_xact_id( T35 ),
       .io_in_1_bits_manager_xact_id( T34 ),
       .io_in_1_bits_is_builtin_type( T33 ),
       .io_in_1_bits_g_type( T32 ),
       .io_in_1_bits_data( T31 ),
       //.io_in_1_bits_client_id(  )
       .io_in_0_ready( gnt_arb_io_in_0_ready ),
       .io_in_0_valid( io_nasti_r_valid ),
       .io_in_0_bits_addr_beat( T22 ),
       .io_in_0_bits_client_xact_id( T21 ),
       .io_in_0_bits_manager_xact_id( T20 ),
       .io_in_0_bits_is_builtin_type( T19 ),
       .io_in_0_bits_g_type( T17 ),
       .io_in_0_bits_data( T14 ),
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_tl_grant_ready ),
       .io_out_valid( gnt_arb_io_out_valid ),
       .io_out_bits_addr_beat( gnt_arb_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( gnt_arb_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( gnt_arb_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( gnt_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( gnt_arb_io_out_bits_g_type ),
       .io_out_bits_data( gnt_arb_io_out_bits_data )
       //.io_out_bits_client_id(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign gnt_arb.io_in_1_bits_client_id = {1{$random}};
    assign gnt_arb.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T10 <= 1'b1;
  if(!T11 && T10 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "NASTI tag error");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T5 <= 1'b1;
  if(!T6 && T5 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "NASTI read error");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "NASTI write error");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else if(T26) begin
      tl_cnt_in <= T25;
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else if(T42) begin
      nasti_cnt_out <= T41;
    end
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else if(T113) begin
      tl_cnt_out <= T112;
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else if(T124) begin
      w_inflight <= 1'h0;
    end else if(T120) begin
      w_inflight <= 1'h1;
    end
  end
endmodule

module ClientTileLinkIOWrapper_1(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [3:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[3:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[3:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[3:0] io_out_release_bits_client_xact_id
    //output io_out_release_bits_voluntary
    //output[2:0] io_out_release_bits_r_type
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module ClientTileLinkEnqueuer(
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [3:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_client_xact_id,
    output io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [3:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [127:0] io_inner_release_bits_data,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[3:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data,
    output io_outer_probe_ready,
    input  io_outer_probe_valid,
    input [25:0] io_outer_probe_bits_addr_block,
    input [1:0] io_outer_probe_bits_p_type,
    input  io_outer_release_ready,
    output io_outer_release_valid,
    output[1:0] io_outer_release_bits_addr_beat,
    output[25:0] io_outer_release_bits_addr_block,
    output[3:0] io_outer_release_bits_client_xact_id,
    output io_outer_release_bits_voluntary,
    output[2:0] io_outer_release_bits_r_type,
    output[127:0] io_outer_release_bits_data
);



  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_acquire_ready = io_outer_acquire_ready;
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [7:0] io_enq_bits_strb,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[7:0] io_deq_bits_strb,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T23;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T24;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire T10;
  wire[73:0] T11;
  reg [73:0] ram [7:0];
  wire[73:0] T12;
  wire[73:0] T13;
  wire[73:0] T14;
  wire[8:0] T15;
  wire[64:0] T16;
  wire[7:0] T17;
  wire T18;
  wire[63:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_strb, io_enq_bits_user};
  assign T16 = {io_enq_bits_data, io_enq_bits_last};
  assign io_deq_bits_strb = T17;
  assign T17 = T11[4'h8:1'h1];
  assign io_deq_bits_last = T18;
  assign T18 = T11[4'h9];
  assign io_deq_bits_data = T19;
  assign T19 = T11[7'h49:4'ha];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [5:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[5:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T25;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T26;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T27;
  wire T8;
  wire T9;
  wire T10;
  wire[73:0] T11;
  reg [73:0] ram [7:0];
  wire[73:0] T12;
  wire[73:0] T13;
  wire[73:0] T14;
  wire[7:0] T15;
  wire[6:0] T16;
  wire[65:0] T17;
  wire[5:0] T18;
  wire T19;
  wire[63:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;
  wire T24;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T25 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T26 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T27 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T17, T15};
  assign T15 = {io_enq_bits_last, T16};
  assign T16 = {io_enq_bits_id, io_enq_bits_user};
  assign T17 = {io_enq_bits_resp, io_enq_bits_data};
  assign io_deq_bits_id = T18;
  assign T18 = T11[3'h6:1'h1];
  assign io_deq_bits_last = T19;
  assign T19 = T11[3'h7];
  assign io_deq_bits_data = T20;
  assign T20 = T11[7'h47:4'h8];
  assign io_deq_bits_resp = T21;
  assign T21 = T11[7'h49:7'h48];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = ptr_match & T23;
  assign T23 = maybe_full ^ 1'h1;
  assign io_enq_ready = T24;
  assign T24 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [5:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[5:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[8:0] T11;
  reg [8:0] ram [1:0];
  wire[8:0] T12;
  wire[8:0] T13;
  wire[8:0] T14;
  wire[6:0] T15;
  wire[5:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_resp, T15};
  assign T15 = {io_enq_bits_id, io_enq_bits_user};
  assign io_deq_bits_id = T16;
  assign T16 = T11[3'h6:1'h1];
  assign io_deq_bits_resp = T17;
  assign T17 = T11[4'h8:3'h7];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module RTC(input clk, input reset,
    input  io_aw_ready,
    output io_aw_valid,
    output[31:0] io_aw_bits_addr,
    output[7:0] io_aw_bits_len,
    output[2:0] io_aw_bits_size,
    output[1:0] io_aw_bits_burst,
    output io_aw_bits_lock,
    output[3:0] io_aw_bits_cache,
    output[2:0] io_aw_bits_prot,
    output[3:0] io_aw_bits_qos,
    output[3:0] io_aw_bits_region,
    output[5:0] io_aw_bits_id,
    output io_aw_bits_user,
    input  io_w_ready,
    output io_w_valid,
    output[63:0] io_w_bits_data,
    output io_w_bits_last,
    output[7:0] io_w_bits_strb,
    output io_w_bits_user,
    output io_b_ready,
    input  io_b_valid,
    input [1:0] io_b_bits_resp,
    input [5:0] io_b_bits_id,
    input  io_b_bits_user,
    input  io_ar_ready,
    output io_ar_valid,
    //output[31:0] io_ar_bits_addr
    //output[7:0] io_ar_bits_len
    //output[2:0] io_ar_bits_size
    //output[1:0] io_ar_bits_burst
    //output io_ar_bits_lock
    //output[3:0] io_ar_bits_cache
    //output[2:0] io_ar_bits_prot
    //output[3:0] io_ar_bits_qos
    //output[3:0] io_ar_bits_region
    //output[5:0] io_ar_bits_id
    //output io_ar_bits_user
    output io_r_ready,
    input  io_r_valid,
    input [1:0] io_r_bits_resp,
    input [63:0] io_r_bits_data,
    input  io_r_bits_last,
    input [5:0] io_r_bits_id,
    input  io_r_bits_user
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  T5;
  wire T6;
  wire T7;
  reg  send_acked_0;
  wire T44;
  wire T8;
  wire T9;
  wire rtc_tick;
  reg [6:0] R10;
  wire[6:0] T45;
  wire[6:0] T11;
  wire[6:0] T12;
  wire T13;
  wire T14;
  wire[1:0] T15;
  wire T16;
  wire T46;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire T21;
  wire[63:0] T22;
  reg [63:0] rtc;
  wire[63:0] T47;
  wire[63:0] T23;
  wire[63:0] T24;
  reg  sending_data;
  wire T48;
  wire T25;
  wire T26;
  wire[5:0] T27;
  wire[5:0] T49;
  wire coreId;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[2:0] T30;
  wire[3:0] T31;
  wire T32;
  wire[1:0] T33;
  wire[2:0] T34;
  wire[7:0] T35;
  wire[31:0] T36;
  wire[31:0] T50;
  reg [30:0] T37;
  reg  sending_addr;
  wire T51;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T5 = 1'b0;
    send_acked_0 = {1{$random}};
    R10 = {1{$random}};
    rtc = {2{$random}};
    sending_data = {1{$random}};
    sending_addr = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_ar_bits_user = {1{$random}};
//  assign io_ar_bits_id = {1{$random}};
//  assign io_ar_bits_region = {1{$random}};
//  assign io_ar_bits_qos = {1{$random}};
//  assign io_ar_bits_prot = {1{$random}};
//  assign io_ar_bits_cache = {1{$random}};
//  assign io_ar_bits_lock = {1{$random}};
//  assign io_ar_bits_burst = {1{$random}};
//  assign io_ar_bits_size = {1{$random}};
//  assign io_ar_bits_len = {1{$random}};
//  assign io_ar_bits_addr = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = io_b_bits_resp == 2'h0;
  assign T4 = io_b_valid ^ 1'h1;
  assign T6 = T7 | reset;
  assign T7 = T18 | send_acked_0;
  assign T44 = reset ? 1'h1 : T8;
  assign T8 = T13 ? 1'h1 : T9;
  assign T9 = rtc_tick ? 1'h0 : send_acked_0;
  assign rtc_tick = R10 == 7'h63;
  assign T45 = reset ? 7'h0 : T11;
  assign T11 = rtc_tick ? 7'h0 : T12;
  assign T12 = R10 + 7'h1;
  assign T13 = T17 & T14;
  assign T14 = T15[1'h0];
  assign T15 = 1'h1 << T16;
  assign T16 = T46;
  assign T46 = io_b_bits_id[1'h0];
  assign T17 = io_b_ready & io_b_valid;
  assign T18 = rtc_tick ^ 1'h1;
  assign io_r_ready = 1'h0;
  assign io_ar_valid = 1'h0;
  assign io_b_ready = 1'h1;
  assign io_w_bits_user = T19;
  assign T19 = 1'h0;
  assign io_w_bits_strb = T20;
  assign T20 = 8'hff;
  assign io_w_bits_last = T21;
  assign T21 = 1'h1;
  assign io_w_bits_data = T22;
  assign T22 = rtc;
  assign T47 = reset ? 64'h0 : T23;
  assign T23 = rtc_tick ? T24 : rtc;
  assign T24 = rtc + 64'h1;
  assign io_w_valid = sending_data;
  assign T48 = reset ? 1'h0 : T25;
  assign T25 = rtc_tick ? 1'h1 : sending_data;
  assign io_aw_bits_user = T26;
  assign T26 = 1'h0;
  assign io_aw_bits_id = T27;
  assign T27 = T49;
  assign T49 = {5'h0, coreId};
  assign coreId = 1'h0;
  assign io_aw_bits_region = T28;
  assign T28 = 4'h0;
  assign io_aw_bits_qos = T29;
  assign T29 = 4'h0;
  assign io_aw_bits_prot = T30;
  assign T30 = 3'h0;
  assign io_aw_bits_cache = T31;
  assign T31 = 4'h0;
  assign io_aw_bits_lock = T32;
  assign T32 = 1'h0;
  assign io_aw_bits_burst = T33;
  assign T33 = 2'h1;
  assign io_aw_bits_size = T34;
  assign T34 = 3'h3;
  assign io_aw_bits_len = T35;
  assign T35 = 8'h0;
  assign io_aw_bits_addr = T36;
  assign T36 = T50;
  assign T50 = {1'h0, T37};
  always @(*) case (coreId)
    0: T37 = 31'h4000b808;
    default: begin
      T37 = 31'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T37 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign io_aw_valid = sending_addr;
  assign T51 = reset ? 1'h0 : T39;
  assign T39 = T43 ? 1'h0 : T40;
  assign T40 = T42 ? 1'h0 : T41;
  assign T41 = rtc_tick ? 1'h1 : sending_addr;
  assign T42 = io_aw_ready & io_aw_valid;
  assign T43 = io_w_ready & io_w_valid;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T5 <= 1'b1;
  if(!T6 && T5 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Not all clocks were updated for rtc tick");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "RTC received NASTI error response");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      send_acked_0 <= 1'h1;
    end else if(T13) begin
      send_acked_0 <= 1'h1;
    end else if(rtc_tick) begin
      send_acked_0 <= 1'h0;
    end
    if(reset) begin
      R10 <= 7'h0;
    end else if(rtc_tick) begin
      R10 <= 7'h0;
    end else begin
      R10 <= T12;
    end
    if(reset) begin
      rtc <= 64'h0;
    end else if(rtc_tick) begin
      rtc <= T24;
    end
    if(reset) begin
      sending_data <= 1'h0;
    end else if(rtc_tick) begin
      sending_data <= 1'h1;
    end
    if(reset) begin
      sending_addr <= 1'h0;
    end else if(T43) begin
      sending_addr <= 1'h0;
    end else if(T42) begin
      sending_addr <= 1'h0;
    end else if(rtc_tick) begin
      sending_addr <= 1'h1;
    end
  end
endmodule

module SmiIONastiReadIOConverter_0(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [5:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[5:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [11:0] addr;
  wire[11:0] T22;
  wire[11:0] T23;
  wire[11:0] T24;
  wire[11:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[5:0] T37;
  reg [5:0] id;
  wire[5:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'he:2'h3];
  assign T25 = addr + 12'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SmiIONastiWriteIOConverter_0(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [5:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[5:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [11:0] addr;
  wire[11:0] T39;
  wire[11:0] T40;
  wire[11:0] T41;
  wire[11:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[5:0] T46;
  reg [5:0] id;
  wire[5:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'he:2'h3];
  assign T42 = addr + 12'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= Smi size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [11:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [11:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[11:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[11:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SmiArbiter_0(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [11:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [11:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[11:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[11:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_1 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SmiIONastiIOConverter_0(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [5:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[5:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [5:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[5:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[5:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[11:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[5:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[11:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[11:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SmiIONastiReadIOConverter_0 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SmiIONastiWriteIOConverter_0 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SmiArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module SmiIONastiReadIOConverter_1(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [5:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[5:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [5:0] addr;
  wire[5:0] T22;
  wire[5:0] T23;
  wire[5:0] T24;
  wire[5:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[5:0] T37;
  reg [5:0] id;
  wire[5:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'h8:2'h3];
  assign T25 = addr + 6'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SmiIONastiWriteIOConverter_1(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [5:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[5:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [5:0] addr;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[5:0] T46;
  reg [5:0] id;
  wire[5:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'h8:2'h3];
  assign T42 = addr + 6'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= Smi size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [5:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [5:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[5:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[5:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SmiArbiter_1(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [5:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [5:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[5:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[5:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_2 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SmiIONastiIOConverter_1(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [5:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[5:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [5:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[5:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[5:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[5:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[5:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[5:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[5:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SmiIONastiReadIOConverter_1 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SmiIONastiWriteIOConverter_1 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SmiArbiter_1 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [5:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[5:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [5:0] io_tiles_cached_0_release_bits_client_xact_id,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [5:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[5:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_uncached_acquire_ready,
    input  io_htif_uncached_acquire_valid,
    input [25:0] io_htif_uncached_acquire_bits_addr_block,
    input [5:0] io_htif_uncached_acquire_bits_client_xact_id,
    input [1:0] io_htif_uncached_acquire_bits_addr_beat,
    input  io_htif_uncached_acquire_bits_is_builtin_type,
    input [2:0] io_htif_uncached_acquire_bits_a_type,
    input [16:0] io_htif_uncached_acquire_bits_union,
    input [127:0] io_htif_uncached_acquire_bits_data,
    input  io_htif_uncached_grant_ready,
    output io_htif_uncached_grant_valid,
    output[1:0] io_htif_uncached_grant_bits_addr_beat,
    output[5:0] io_htif_uncached_grant_bits_client_xact_id,
    output[3:0] io_htif_uncached_grant_bits_manager_xact_id,
    output io_htif_uncached_grant_bits_is_builtin_type,
    output[3:0] io_htif_uncached_grant_bits_g_type,
    output[127:0] io_htif_uncached_grant_bits_data,
    input  io_incoherent_0,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[5:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [5:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[5:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [5:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    input  io_mem_backup_req_ready,
    output io_mem_backup_req_valid,
    output[15:0] io_mem_backup_req_bits,
    input  io_mem_backup_resp_valid,
    input [15:0] io_mem_backup_resp_bits,
    input  io_mem_backup_en,
    input  io_memory_channel_mux_select,
    input  io_csr_0_req_ready,
    output io_csr_0_req_valid,
    output io_csr_0_req_bits_rw,
    output[11:0] io_csr_0_req_bits_addr,
    output[63:0] io_csr_0_req_bits_data,
    output io_csr_0_resp_ready,
    input  io_csr_0_resp_valid,
    input [63:0] io_csr_0_resp_bits,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits,
    input  io_deviceTree_aw_ready,
    output io_deviceTree_aw_valid,
    output[31:0] io_deviceTree_aw_bits_addr,
    output[7:0] io_deviceTree_aw_bits_len,
    output[2:0] io_deviceTree_aw_bits_size,
    output[1:0] io_deviceTree_aw_bits_burst,
    output io_deviceTree_aw_bits_lock,
    output[3:0] io_deviceTree_aw_bits_cache,
    output[2:0] io_deviceTree_aw_bits_prot,
    output[3:0] io_deviceTree_aw_bits_qos,
    output[3:0] io_deviceTree_aw_bits_region,
    output[5:0] io_deviceTree_aw_bits_id,
    output io_deviceTree_aw_bits_user,
    input  io_deviceTree_w_ready,
    output io_deviceTree_w_valid,
    output[63:0] io_deviceTree_w_bits_data,
    output io_deviceTree_w_bits_last,
    output[7:0] io_deviceTree_w_bits_strb,
    output io_deviceTree_w_bits_user,
    output io_deviceTree_b_ready,
    input  io_deviceTree_b_valid,
    input [1:0] io_deviceTree_b_bits_resp,
    input [5:0] io_deviceTree_b_bits_id,
    input  io_deviceTree_b_bits_user,
    input  io_deviceTree_ar_ready,
    output io_deviceTree_ar_valid,
    output[31:0] io_deviceTree_ar_bits_addr,
    output[7:0] io_deviceTree_ar_bits_len,
    output[2:0] io_deviceTree_ar_bits_size,
    output[1:0] io_deviceTree_ar_bits_burst,
    output io_deviceTree_ar_bits_lock,
    output[3:0] io_deviceTree_ar_bits_cache,
    output[2:0] io_deviceTree_ar_bits_prot,
    output[3:0] io_deviceTree_ar_bits_qos,
    output[3:0] io_deviceTree_ar_bits_region,
    output[5:0] io_deviceTree_ar_bits_id,
    output io_deviceTree_ar_bits_user,
    output io_deviceTree_r_ready,
    input  io_deviceTree_r_valid,
    input [1:0] io_deviceTree_r_bits_resp,
    input [63:0] io_deviceTree_r_bits_data,
    input  io_deviceTree_r_bits_last,
    input [5:0] io_deviceTree_r_bits_id,
    input  io_deviceTree_r_bits_user
);

  wire ClientTileLinkIOWrapper_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block;
  wire[5:0] ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_io_out_release_valid;
  wire ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_1_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block;
  wire[5:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_1_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_1_io_out_release_valid;
  wire mmioManager_io_inner_acquire_ready;
  wire mmioManager_io_inner_grant_valid;
  wire[1:0] mmioManager_io_inner_grant_bits_addr_beat;
  wire[5:0] mmioManager_io_inner_grant_bits_client_xact_id;
  wire[3:0] mmioManager_io_inner_grant_bits_manager_xact_id;
  wire mmioManager_io_inner_grant_bits_is_builtin_type;
  wire[3:0] mmioManager_io_inner_grant_bits_g_type;
  wire[127:0] mmioManager_io_inner_grant_bits_data;
  wire[1:0] mmioManager_io_inner_grant_bits_client_id;
  wire mmioManager_io_inner_finish_ready;
  wire mmioManager_io_inner_probe_valid;
  wire mmioManager_io_inner_release_ready;
  wire mmioManager_io_outer_acquire_valid;
  wire[25:0] mmioManager_io_outer_acquire_bits_addr_block;
  wire[3:0] mmioManager_io_outer_acquire_bits_client_xact_id;
  wire[1:0] mmioManager_io_outer_acquire_bits_addr_beat;
  wire mmioManager_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] mmioManager_io_outer_acquire_bits_a_type;
  wire[16:0] mmioManager_io_outer_acquire_bits_union;
  wire[127:0] mmioManager_io_outer_acquire_bits_data;
  wire mmioManager_io_outer_grant_ready;
  wire ClientTileLinkIOWrapper_2_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_2_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block;
  wire[3:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_2_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_2_io_out_release_valid;
  wire ClientTileLinkEnqueuer_io_inner_acquire_ready;
  wire ClientTileLinkEnqueuer_io_inner_grant_valid;
  wire[1:0] ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat;
  wire[3:0] ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id;
  wire ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id;
  wire ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkEnqueuer_io_inner_grant_bits_g_type;
  wire[127:0] ClientTileLinkEnqueuer_io_inner_grant_bits_data;
  wire ClientTileLinkEnqueuer_io_inner_probe_valid;
  wire[25:0] ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block;
  wire[1:0] ClientTileLinkEnqueuer_io_inner_probe_bits_p_type;
  wire ClientTileLinkEnqueuer_io_inner_release_ready;
  wire ClientTileLinkEnqueuer_io_outer_acquire_valid;
  wire[25:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block;
  wire[3:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat;
  wire ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type;
  wire[16:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_union;
  wire[127:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_data;
  wire ClientTileLinkEnqueuer_io_outer_grant_ready;
  wire ClientTileLinkEnqueuer_io_outer_probe_ready;
  wire ClientTileLinkEnqueuer_io_outer_release_valid;
  wire[1:0] ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat;
  wire[25:0] ClientTileLinkEnqueuer_io_outer_release_bits_addr_block;
  wire[3:0] ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id;
  wire ClientTileLinkEnqueuer_io_outer_release_bits_voluntary;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_release_bits_r_type;
  wire[127:0] ClientTileLinkEnqueuer_io_outer_release_bits_data;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[31:0] Queue_io_deq_bits_addr;
  wire[7:0] Queue_io_deq_bits_len;
  wire[2:0] Queue_io_deq_bits_size;
  wire[1:0] Queue_io_deq_bits_burst;
  wire Queue_io_deq_bits_lock;
  wire[3:0] Queue_io_deq_bits_cache;
  wire[2:0] Queue_io_deq_bits_prot;
  wire[3:0] Queue_io_deq_bits_qos;
  wire[3:0] Queue_io_deq_bits_region;
  wire[5:0] Queue_io_deq_bits_id;
  wire Queue_io_deq_bits_user;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[31:0] Queue_1_io_deq_bits_addr;
  wire[7:0] Queue_1_io_deq_bits_len;
  wire[2:0] Queue_1_io_deq_bits_size;
  wire[1:0] Queue_1_io_deq_bits_burst;
  wire Queue_1_io_deq_bits_lock;
  wire[3:0] Queue_1_io_deq_bits_cache;
  wire[2:0] Queue_1_io_deq_bits_prot;
  wire[3:0] Queue_1_io_deq_bits_qos;
  wire[3:0] Queue_1_io_deq_bits_region;
  wire[5:0] Queue_1_io_deq_bits_id;
  wire Queue_1_io_deq_bits_user;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[63:0] Queue_2_io_deq_bits_data;
  wire Queue_2_io_deq_bits_last;
  wire[7:0] Queue_2_io_deq_bits_strb;
  wire Queue_2_io_deq_bits_user;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_resp;
  wire[63:0] Queue_3_io_deq_bits_data;
  wire Queue_3_io_deq_bits_last;
  wire[5:0] Queue_3_io_deq_bits_id;
  wire Queue_3_io_deq_bits_user;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_resp;
  wire[5:0] Queue_4_io_deq_bits_id;
  wire Queue_4_io_deq_bits_user;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[31:0] Queue_5_io_deq_bits_addr;
  wire[7:0] Queue_5_io_deq_bits_len;
  wire[2:0] Queue_5_io_deq_bits_size;
  wire[1:0] Queue_5_io_deq_bits_burst;
  wire Queue_5_io_deq_bits_lock;
  wire[3:0] Queue_5_io_deq_bits_cache;
  wire[2:0] Queue_5_io_deq_bits_prot;
  wire[3:0] Queue_5_io_deq_bits_qos;
  wire[3:0] Queue_5_io_deq_bits_region;
  wire[5:0] Queue_5_io_deq_bits_id;
  wire Queue_5_io_deq_bits_user;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[31:0] Queue_6_io_deq_bits_addr;
  wire[7:0] Queue_6_io_deq_bits_len;
  wire[2:0] Queue_6_io_deq_bits_size;
  wire[1:0] Queue_6_io_deq_bits_burst;
  wire Queue_6_io_deq_bits_lock;
  wire[3:0] Queue_6_io_deq_bits_cache;
  wire[2:0] Queue_6_io_deq_bits_prot;
  wire[3:0] Queue_6_io_deq_bits_qos;
  wire[3:0] Queue_6_io_deq_bits_region;
  wire[5:0] Queue_6_io_deq_bits_id;
  wire Queue_6_io_deq_bits_user;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[63:0] Queue_7_io_deq_bits_data;
  wire Queue_7_io_deq_bits_last;
  wire[7:0] Queue_7_io_deq_bits_strb;
  wire Queue_7_io_deq_bits_user;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_resp;
  wire[63:0] Queue_8_io_deq_bits_data;
  wire Queue_8_io_deq_bits_last;
  wire[5:0] Queue_8_io_deq_bits_id;
  wire Queue_8_io_deq_bits_user;
  wire Queue_9_io_enq_ready;
  wire Queue_9_io_deq_valid;
  wire[1:0] Queue_9_io_deq_bits_resp;
  wire[5:0] Queue_9_io_deq_bits_id;
  wire Queue_9_io_deq_bits_user;
  wire rtc_io_aw_valid;
  wire[31:0] rtc_io_aw_bits_addr;
  wire[7:0] rtc_io_aw_bits_len;
  wire[2:0] rtc_io_aw_bits_size;
  wire[1:0] rtc_io_aw_bits_burst;
  wire rtc_io_aw_bits_lock;
  wire[3:0] rtc_io_aw_bits_cache;
  wire[2:0] rtc_io_aw_bits_prot;
  wire[3:0] rtc_io_aw_bits_qos;
  wire[3:0] rtc_io_aw_bits_region;
  wire[5:0] rtc_io_aw_bits_id;
  wire rtc_io_aw_bits_user;
  wire rtc_io_w_valid;
  wire[63:0] rtc_io_w_bits_data;
  wire rtc_io_w_bits_last;
  wire[7:0] rtc_io_w_bits_strb;
  wire rtc_io_w_bits_user;
  wire rtc_io_b_ready;
  wire rtc_io_ar_valid;
  wire rtc_io_r_ready;
  wire mem_ic_io_masters_0_aw_ready;
  wire mem_ic_io_masters_0_w_ready;
  wire mem_ic_io_masters_0_b_valid;
  wire[1:0] mem_ic_io_masters_0_b_bits_resp;
  wire[5:0] mem_ic_io_masters_0_b_bits_id;
  wire mem_ic_io_masters_0_b_bits_user;
  wire mem_ic_io_masters_0_ar_ready;
  wire mem_ic_io_masters_0_r_valid;
  wire[1:0] mem_ic_io_masters_0_r_bits_resp;
  wire[63:0] mem_ic_io_masters_0_r_bits_data;
  wire mem_ic_io_masters_0_r_bits_last;
  wire[5:0] mem_ic_io_masters_0_r_bits_id;
  wire mem_ic_io_masters_0_r_bits_user;
  wire mem_ic_io_slaves_0_aw_valid;
  wire[31:0] mem_ic_io_slaves_0_aw_bits_addr;
  wire[7:0] mem_ic_io_slaves_0_aw_bits_len;
  wire[2:0] mem_ic_io_slaves_0_aw_bits_size;
  wire[1:0] mem_ic_io_slaves_0_aw_bits_burst;
  wire mem_ic_io_slaves_0_aw_bits_lock;
  wire[3:0] mem_ic_io_slaves_0_aw_bits_cache;
  wire[2:0] mem_ic_io_slaves_0_aw_bits_prot;
  wire[3:0] mem_ic_io_slaves_0_aw_bits_qos;
  wire[3:0] mem_ic_io_slaves_0_aw_bits_region;
  wire[5:0] mem_ic_io_slaves_0_aw_bits_id;
  wire mem_ic_io_slaves_0_aw_bits_user;
  wire mem_ic_io_slaves_0_w_valid;
  wire[63:0] mem_ic_io_slaves_0_w_bits_data;
  wire mem_ic_io_slaves_0_w_bits_last;
  wire[7:0] mem_ic_io_slaves_0_w_bits_strb;
  wire mem_ic_io_slaves_0_w_bits_user;
  wire mem_ic_io_slaves_0_b_ready;
  wire mem_ic_io_slaves_0_ar_valid;
  wire[31:0] mem_ic_io_slaves_0_ar_bits_addr;
  wire[7:0] mem_ic_io_slaves_0_ar_bits_len;
  wire[2:0] mem_ic_io_slaves_0_ar_bits_size;
  wire[1:0] mem_ic_io_slaves_0_ar_bits_burst;
  wire mem_ic_io_slaves_0_ar_bits_lock;
  wire[3:0] mem_ic_io_slaves_0_ar_bits_cache;
  wire[2:0] mem_ic_io_slaves_0_ar_bits_prot;
  wire[3:0] mem_ic_io_slaves_0_ar_bits_qos;
  wire[3:0] mem_ic_io_slaves_0_ar_bits_region;
  wire[5:0] mem_ic_io_slaves_0_ar_bits_id;
  wire mem_ic_io_slaves_0_ar_bits_user;
  wire mem_ic_io_slaves_0_r_ready;
  wire ClientTileLinkIOUnwrapper_io_in_acquire_ready;
  wire ClientTileLinkIOUnwrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat;
  wire[3:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOUnwrapper_io_in_probe_valid;
  wire ClientTileLinkIOUnwrapper_io_in_release_ready;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block;
  wire[3:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOUnwrapper_io_out_grant_ready;
  wire TileLinkIONarrower_io_in_acquire_ready;
  wire TileLinkIONarrower_io_in_grant_valid;
  wire[1:0] TileLinkIONarrower_io_in_grant_bits_addr_beat;
  wire[3:0] TileLinkIONarrower_io_in_grant_bits_client_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_manager_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_is_builtin_type;
  wire[3:0] TileLinkIONarrower_io_in_grant_bits_g_type;
  wire[127:0] TileLinkIONarrower_io_in_grant_bits_data;
  wire TileLinkIONarrower_io_out_acquire_valid;
  wire[25:0] TileLinkIONarrower_io_out_acquire_bits_addr_block;
  wire[3:0] TileLinkIONarrower_io_out_acquire_bits_client_xact_id;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_addr_beat;
  wire TileLinkIONarrower_io_out_acquire_bits_is_builtin_type;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_a_type;
  wire[11:0] TileLinkIONarrower_io_out_acquire_bits_union;
  wire[63:0] TileLinkIONarrower_io_out_acquire_bits_data;
  wire TileLinkIONarrower_io_out_grant_ready;
  wire NastiIOTileLinkIOConverter_io_tl_acquire_ready;
  wire NastiIOTileLinkIOConverter_io_tl_grant_valid;
  wire[2:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat;
  wire[3:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type;
  wire[3:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type;
  wire[63:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_region;
  wire[5:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_w_valid;
  wire[63:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_last;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_strb;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_b_ready;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_region;
  wire[5:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_r_ready;
  wire mmio_narrow_io_in_acquire_ready;
  wire mmio_narrow_io_in_grant_valid;
  wire[1:0] mmio_narrow_io_in_grant_bits_addr_beat;
  wire[3:0] mmio_narrow_io_in_grant_bits_client_xact_id;
  wire mmio_narrow_io_in_grant_bits_manager_xact_id;
  wire mmio_narrow_io_in_grant_bits_is_builtin_type;
  wire[3:0] mmio_narrow_io_in_grant_bits_g_type;
  wire[127:0] mmio_narrow_io_in_grant_bits_data;
  wire mmio_narrow_io_out_acquire_valid;
  wire[25:0] mmio_narrow_io_out_acquire_bits_addr_block;
  wire[3:0] mmio_narrow_io_out_acquire_bits_client_xact_id;
  wire[2:0] mmio_narrow_io_out_acquire_bits_addr_beat;
  wire mmio_narrow_io_out_acquire_bits_is_builtin_type;
  wire[2:0] mmio_narrow_io_out_acquire_bits_a_type;
  wire[11:0] mmio_narrow_io_out_acquire_bits_union;
  wire[63:0] mmio_narrow_io_out_acquire_bits_data;
  wire mmio_narrow_io_out_grant_ready;
  wire mmio_conv_io_tl_acquire_ready;
  wire mmio_conv_io_tl_grant_valid;
  wire[2:0] mmio_conv_io_tl_grant_bits_addr_beat;
  wire[3:0] mmio_conv_io_tl_grant_bits_client_xact_id;
  wire mmio_conv_io_tl_grant_bits_manager_xact_id;
  wire mmio_conv_io_tl_grant_bits_is_builtin_type;
  wire[3:0] mmio_conv_io_tl_grant_bits_g_type;
  wire[63:0] mmio_conv_io_tl_grant_bits_data;
  wire mmio_conv_io_nasti_aw_valid;
  wire[31:0] mmio_conv_io_nasti_aw_bits_addr;
  wire[7:0] mmio_conv_io_nasti_aw_bits_len;
  wire[2:0] mmio_conv_io_nasti_aw_bits_size;
  wire[1:0] mmio_conv_io_nasti_aw_bits_burst;
  wire mmio_conv_io_nasti_aw_bits_lock;
  wire[3:0] mmio_conv_io_nasti_aw_bits_cache;
  wire[2:0] mmio_conv_io_nasti_aw_bits_prot;
  wire[3:0] mmio_conv_io_nasti_aw_bits_qos;
  wire[3:0] mmio_conv_io_nasti_aw_bits_region;
  wire[5:0] mmio_conv_io_nasti_aw_bits_id;
  wire mmio_conv_io_nasti_aw_bits_user;
  wire mmio_conv_io_nasti_w_valid;
  wire[63:0] mmio_conv_io_nasti_w_bits_data;
  wire mmio_conv_io_nasti_w_bits_last;
  wire[7:0] mmio_conv_io_nasti_w_bits_strb;
  wire mmio_conv_io_nasti_w_bits_user;
  wire mmio_conv_io_nasti_b_ready;
  wire mmio_conv_io_nasti_ar_valid;
  wire[31:0] mmio_conv_io_nasti_ar_bits_addr;
  wire[7:0] mmio_conv_io_nasti_ar_bits_len;
  wire[2:0] mmio_conv_io_nasti_ar_bits_size;
  wire[1:0] mmio_conv_io_nasti_ar_bits_burst;
  wire mmio_conv_io_nasti_ar_bits_lock;
  wire[3:0] mmio_conv_io_nasti_ar_bits_cache;
  wire[2:0] mmio_conv_io_nasti_ar_bits_prot;
  wire[3:0] mmio_conv_io_nasti_ar_bits_qos;
  wire[3:0] mmio_conv_io_nasti_ar_bits_region;
  wire[5:0] mmio_conv_io_nasti_ar_bits_id;
  wire mmio_conv_io_nasti_ar_bits_user;
  wire mmio_conv_io_nasti_r_ready;
  wire L2BroadcastHub_io_inner_acquire_ready;
  wire L2BroadcastHub_io_inner_grant_valid;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_addr_beat;
  wire[5:0] L2BroadcastHub_io_inner_grant_bits_client_xact_id;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_manager_xact_id;
  wire L2BroadcastHub_io_inner_grant_bits_is_builtin_type;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_g_type;
  wire[127:0] L2BroadcastHub_io_inner_grant_bits_data;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_id;
  wire L2BroadcastHub_io_inner_finish_ready;
  wire L2BroadcastHub_io_inner_probe_valid;
  wire[25:0] L2BroadcastHub_io_inner_probe_bits_addr_block;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_p_type;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_client_id;
  wire L2BroadcastHub_io_inner_release_ready;
  wire L2BroadcastHub_io_outer_acquire_valid;
  wire[25:0] L2BroadcastHub_io_outer_acquire_bits_addr_block;
  wire[3:0] L2BroadcastHub_io_outer_acquire_bits_client_xact_id;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_addr_beat;
  wire L2BroadcastHub_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_a_type;
  wire[16:0] L2BroadcastHub_io_outer_acquire_bits_union;
  wire[127:0] L2BroadcastHub_io_outer_acquire_bits_data;
  wire L2BroadcastHub_io_outer_grant_ready;
  wire SmiIONastiIOConverter_io_nasti_aw_ready;
  wire SmiIONastiIOConverter_io_nasti_w_ready;
  wire SmiIONastiIOConverter_io_nasti_b_valid;
  wire[1:0] SmiIONastiIOConverter_io_nasti_b_bits_resp;
  wire[5:0] SmiIONastiIOConverter_io_nasti_b_bits_id;
  wire SmiIONastiIOConverter_io_nasti_b_bits_user;
  wire SmiIONastiIOConverter_io_nasti_ar_ready;
  wire SmiIONastiIOConverter_io_nasti_r_valid;
  wire[1:0] SmiIONastiIOConverter_io_nasti_r_bits_resp;
  wire[63:0] SmiIONastiIOConverter_io_nasti_r_bits_data;
  wire SmiIONastiIOConverter_io_nasti_r_bits_last;
  wire[5:0] SmiIONastiIOConverter_io_nasti_r_bits_id;
  wire SmiIONastiIOConverter_io_nasti_r_bits_user;
  wire SmiIONastiIOConverter_io_smi_req_valid;
  wire SmiIONastiIOConverter_io_smi_req_bits_rw;
  wire[11:0] SmiIONastiIOConverter_io_smi_req_bits_addr;
  wire[63:0] SmiIONastiIOConverter_io_smi_req_bits_data;
  wire SmiIONastiIOConverter_io_smi_resp_ready;
  wire scr_conv_io_nasti_aw_ready;
  wire scr_conv_io_nasti_w_ready;
  wire scr_conv_io_nasti_b_valid;
  wire[1:0] scr_conv_io_nasti_b_bits_resp;
  wire[5:0] scr_conv_io_nasti_b_bits_id;
  wire scr_conv_io_nasti_b_bits_user;
  wire scr_conv_io_nasti_ar_ready;
  wire scr_conv_io_nasti_r_valid;
  wire[1:0] scr_conv_io_nasti_r_bits_resp;
  wire[63:0] scr_conv_io_nasti_r_bits_data;
  wire scr_conv_io_nasti_r_bits_last;
  wire[5:0] scr_conv_io_nasti_r_bits_id;
  wire scr_conv_io_nasti_r_bits_user;
  wire scr_conv_io_smi_req_valid;
  wire scr_conv_io_smi_req_bits_rw;
  wire[5:0] scr_conv_io_smi_req_bits_addr;
  wire[63:0] scr_conv_io_smi_req_bits_data;
  wire scr_conv_io_smi_resp_ready;
  wire l1tol2net_io_clients_2_acquire_ready;
  wire l1tol2net_io_clients_2_grant_valid;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_addr_beat;
  wire[5:0] l1tol2net_io_clients_2_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_2_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_2_grant_bits_data;
  wire l1tol2net_io_clients_2_probe_valid;
  wire[25:0] l1tol2net_io_clients_2_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_2_probe_bits_p_type;
  wire l1tol2net_io_clients_2_release_ready;
  wire l1tol2net_io_clients_1_acquire_ready;
  wire l1tol2net_io_clients_1_grant_valid;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_addr_beat;
  wire[5:0] l1tol2net_io_clients_1_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_1_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_1_grant_bits_data;
  wire l1tol2net_io_clients_1_probe_valid;
  wire[25:0] l1tol2net_io_clients_1_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_1_probe_bits_p_type;
  wire l1tol2net_io_clients_1_release_ready;
  wire l1tol2net_io_clients_0_acquire_ready;
  wire l1tol2net_io_clients_0_grant_valid;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_addr_beat;
  wire[5:0] l1tol2net_io_clients_0_grant_bits_client_xact_id;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_0_grant_bits_data;
  wire l1tol2net_io_clients_0_probe_valid;
  wire[25:0] l1tol2net_io_clients_0_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_0_probe_bits_p_type;
  wire l1tol2net_io_clients_0_release_ready;
  wire l1tol2net_io_managers_1_acquire_valid;
  wire[25:0] l1tol2net_io_managers_1_acquire_bits_addr_block;
  wire[5:0] l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_1_acquire_bits_addr_beat;
  wire l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  wire[2:0] l1tol2net_io_managers_1_acquire_bits_a_type;
  wire[16:0] l1tol2net_io_managers_1_acquire_bits_union;
  wire[127:0] l1tol2net_io_managers_1_acquire_bits_data;
  wire[1:0] l1tol2net_io_managers_1_acquire_bits_client_id;
  wire l1tol2net_io_managers_1_grant_ready;
  wire l1tol2net_io_managers_1_finish_valid;
  wire[3:0] l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  wire l1tol2net_io_managers_1_probe_ready;
  wire l1tol2net_io_managers_1_release_valid;
  wire[1:0] l1tol2net_io_managers_1_release_bits_addr_beat;
  wire[25:0] l1tol2net_io_managers_1_release_bits_addr_block;
  wire[5:0] l1tol2net_io_managers_1_release_bits_client_xact_id;
  wire l1tol2net_io_managers_1_release_bits_voluntary;
  wire[2:0] l1tol2net_io_managers_1_release_bits_r_type;
  wire[127:0] l1tol2net_io_managers_1_release_bits_data;
  wire[1:0] l1tol2net_io_managers_1_release_bits_client_id;
  wire l1tol2net_io_managers_0_acquire_valid;
  wire[25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire[5:0] l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire[2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire[16:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire[127:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_id;
  wire l1tol2net_io_managers_0_grant_ready;
  wire l1tol2net_io_managers_0_finish_valid;
  wire[3:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire l1tol2net_io_managers_0_probe_ready;
  wire l1tol2net_io_managers_0_release_valid;
  wire[1:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire[25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire[5:0] l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire l1tol2net_io_managers_0_release_bits_voluntary;
  wire[2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire[127:0] l1tol2net_io_managers_0_release_bits_data;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_id;
  wire mmio_ic_io_masters_1_aw_ready;
  wire mmio_ic_io_masters_1_w_ready;
  wire mmio_ic_io_masters_1_b_valid;
  wire[1:0] mmio_ic_io_masters_1_b_bits_resp;
  wire[5:0] mmio_ic_io_masters_1_b_bits_id;
  wire mmio_ic_io_masters_1_b_bits_user;
  wire mmio_ic_io_masters_1_ar_ready;
  wire mmio_ic_io_masters_1_r_valid;
  wire[1:0] mmio_ic_io_masters_1_r_bits_resp;
  wire[63:0] mmio_ic_io_masters_1_r_bits_data;
  wire mmio_ic_io_masters_1_r_bits_last;
  wire[5:0] mmio_ic_io_masters_1_r_bits_id;
  wire mmio_ic_io_masters_1_r_bits_user;
  wire mmio_ic_io_masters_0_aw_ready;
  wire mmio_ic_io_masters_0_w_ready;
  wire mmio_ic_io_masters_0_b_valid;
  wire[1:0] mmio_ic_io_masters_0_b_bits_resp;
  wire[5:0] mmio_ic_io_masters_0_b_bits_id;
  wire mmio_ic_io_masters_0_b_bits_user;
  wire mmio_ic_io_masters_0_ar_ready;
  wire mmio_ic_io_masters_0_r_valid;
  wire[1:0] mmio_ic_io_masters_0_r_bits_resp;
  wire[63:0] mmio_ic_io_masters_0_r_bits_data;
  wire mmio_ic_io_masters_0_r_bits_last;
  wire[5:0] mmio_ic_io_masters_0_r_bits_id;
  wire mmio_ic_io_masters_0_r_bits_user;
  wire mmio_ic_io_slaves_2_aw_valid;
  wire[31:0] mmio_ic_io_slaves_2_aw_bits_addr;
  wire[7:0] mmio_ic_io_slaves_2_aw_bits_len;
  wire[2:0] mmio_ic_io_slaves_2_aw_bits_size;
  wire[1:0] mmio_ic_io_slaves_2_aw_bits_burst;
  wire mmio_ic_io_slaves_2_aw_bits_lock;
  wire[3:0] mmio_ic_io_slaves_2_aw_bits_cache;
  wire[2:0] mmio_ic_io_slaves_2_aw_bits_prot;
  wire[3:0] mmio_ic_io_slaves_2_aw_bits_qos;
  wire[3:0] mmio_ic_io_slaves_2_aw_bits_region;
  wire[5:0] mmio_ic_io_slaves_2_aw_bits_id;
  wire mmio_ic_io_slaves_2_aw_bits_user;
  wire mmio_ic_io_slaves_2_w_valid;
  wire[63:0] mmio_ic_io_slaves_2_w_bits_data;
  wire mmio_ic_io_slaves_2_w_bits_last;
  wire[7:0] mmio_ic_io_slaves_2_w_bits_strb;
  wire mmio_ic_io_slaves_2_w_bits_user;
  wire mmio_ic_io_slaves_2_b_ready;
  wire mmio_ic_io_slaves_2_ar_valid;
  wire[31:0] mmio_ic_io_slaves_2_ar_bits_addr;
  wire[7:0] mmio_ic_io_slaves_2_ar_bits_len;
  wire[2:0] mmio_ic_io_slaves_2_ar_bits_size;
  wire[1:0] mmio_ic_io_slaves_2_ar_bits_burst;
  wire mmio_ic_io_slaves_2_ar_bits_lock;
  wire[3:0] mmio_ic_io_slaves_2_ar_bits_cache;
  wire[2:0] mmio_ic_io_slaves_2_ar_bits_prot;
  wire[3:0] mmio_ic_io_slaves_2_ar_bits_qos;
  wire[3:0] mmio_ic_io_slaves_2_ar_bits_region;
  wire[5:0] mmio_ic_io_slaves_2_ar_bits_id;
  wire mmio_ic_io_slaves_2_ar_bits_user;
  wire mmio_ic_io_slaves_2_r_ready;
  wire mmio_ic_io_slaves_1_aw_valid;
  wire[31:0] mmio_ic_io_slaves_1_aw_bits_addr;
  wire[7:0] mmio_ic_io_slaves_1_aw_bits_len;
  wire[2:0] mmio_ic_io_slaves_1_aw_bits_size;
  wire[1:0] mmio_ic_io_slaves_1_aw_bits_burst;
  wire mmio_ic_io_slaves_1_aw_bits_lock;
  wire[3:0] mmio_ic_io_slaves_1_aw_bits_cache;
  wire[2:0] mmio_ic_io_slaves_1_aw_bits_prot;
  wire[3:0] mmio_ic_io_slaves_1_aw_bits_qos;
  wire[3:0] mmio_ic_io_slaves_1_aw_bits_region;
  wire[5:0] mmio_ic_io_slaves_1_aw_bits_id;
  wire mmio_ic_io_slaves_1_aw_bits_user;
  wire mmio_ic_io_slaves_1_w_valid;
  wire[63:0] mmio_ic_io_slaves_1_w_bits_data;
  wire mmio_ic_io_slaves_1_w_bits_last;
  wire[7:0] mmio_ic_io_slaves_1_w_bits_strb;
  wire mmio_ic_io_slaves_1_w_bits_user;
  wire mmio_ic_io_slaves_1_b_ready;
  wire mmio_ic_io_slaves_1_ar_valid;
  wire[31:0] mmio_ic_io_slaves_1_ar_bits_addr;
  wire[7:0] mmio_ic_io_slaves_1_ar_bits_len;
  wire[2:0] mmio_ic_io_slaves_1_ar_bits_size;
  wire[1:0] mmio_ic_io_slaves_1_ar_bits_burst;
  wire mmio_ic_io_slaves_1_ar_bits_lock;
  wire[3:0] mmio_ic_io_slaves_1_ar_bits_cache;
  wire[2:0] mmio_ic_io_slaves_1_ar_bits_prot;
  wire[3:0] mmio_ic_io_slaves_1_ar_bits_qos;
  wire[3:0] mmio_ic_io_slaves_1_ar_bits_region;
  wire[5:0] mmio_ic_io_slaves_1_ar_bits_id;
  wire mmio_ic_io_slaves_1_ar_bits_user;
  wire mmio_ic_io_slaves_1_r_ready;
  wire mmio_ic_io_slaves_0_aw_valid;
  wire[31:0] mmio_ic_io_slaves_0_aw_bits_addr;
  wire[7:0] mmio_ic_io_slaves_0_aw_bits_len;
  wire[2:0] mmio_ic_io_slaves_0_aw_bits_size;
  wire[1:0] mmio_ic_io_slaves_0_aw_bits_burst;
  wire mmio_ic_io_slaves_0_aw_bits_lock;
  wire[3:0] mmio_ic_io_slaves_0_aw_bits_cache;
  wire[2:0] mmio_ic_io_slaves_0_aw_bits_prot;
  wire[3:0] mmio_ic_io_slaves_0_aw_bits_qos;
  wire[3:0] mmio_ic_io_slaves_0_aw_bits_region;
  wire[5:0] mmio_ic_io_slaves_0_aw_bits_id;
  wire mmio_ic_io_slaves_0_aw_bits_user;
  wire mmio_ic_io_slaves_0_w_valid;
  wire[63:0] mmio_ic_io_slaves_0_w_bits_data;
  wire mmio_ic_io_slaves_0_w_bits_last;
  wire[7:0] mmio_ic_io_slaves_0_w_bits_strb;
  wire mmio_ic_io_slaves_0_w_bits_user;
  wire mmio_ic_io_slaves_0_b_ready;
  wire mmio_ic_io_slaves_0_ar_valid;
  wire[31:0] mmio_ic_io_slaves_0_ar_bits_addr;
  wire[7:0] mmio_ic_io_slaves_0_ar_bits_len;
  wire[2:0] mmio_ic_io_slaves_0_ar_bits_size;
  wire[1:0] mmio_ic_io_slaves_0_ar_bits_burst;
  wire mmio_ic_io_slaves_0_ar_bits_lock;
  wire[3:0] mmio_ic_io_slaves_0_ar_bits_cache;
  wire[2:0] mmio_ic_io_slaves_0_ar_bits_prot;
  wire[3:0] mmio_ic_io_slaves_0_ar_bits_qos;
  wire[3:0] mmio_ic_io_slaves_0_ar_bits_region;
  wire[5:0] mmio_ic_io_slaves_0_ar_bits_id;
  wire mmio_ic_io_slaves_0_ar_bits_user;
  wire mmio_ic_io_slaves_0_r_ready;


`ifndef SYNTHESIS
// synthesis translate_off
  assign io_mem_backup_req_bits = {1{$random}};
// synthesis translate_on
`endif
  assign io_deviceTree_r_ready = mmio_ic_io_slaves_0_r_ready;
  assign io_deviceTree_ar_bits_user = mmio_ic_io_slaves_0_ar_bits_user;
  assign io_deviceTree_ar_bits_id = mmio_ic_io_slaves_0_ar_bits_id;
  assign io_deviceTree_ar_bits_region = mmio_ic_io_slaves_0_ar_bits_region;
  assign io_deviceTree_ar_bits_qos = mmio_ic_io_slaves_0_ar_bits_qos;
  assign io_deviceTree_ar_bits_prot = mmio_ic_io_slaves_0_ar_bits_prot;
  assign io_deviceTree_ar_bits_cache = mmio_ic_io_slaves_0_ar_bits_cache;
  assign io_deviceTree_ar_bits_lock = mmio_ic_io_slaves_0_ar_bits_lock;
  assign io_deviceTree_ar_bits_burst = mmio_ic_io_slaves_0_ar_bits_burst;
  assign io_deviceTree_ar_bits_size = mmio_ic_io_slaves_0_ar_bits_size;
  assign io_deviceTree_ar_bits_len = mmio_ic_io_slaves_0_ar_bits_len;
  assign io_deviceTree_ar_bits_addr = mmio_ic_io_slaves_0_ar_bits_addr;
  assign io_deviceTree_ar_valid = mmio_ic_io_slaves_0_ar_valid;
  assign io_deviceTree_b_ready = mmio_ic_io_slaves_0_b_ready;
  assign io_deviceTree_w_bits_user = mmio_ic_io_slaves_0_w_bits_user;
  assign io_deviceTree_w_bits_strb = mmio_ic_io_slaves_0_w_bits_strb;
  assign io_deviceTree_w_bits_last = mmio_ic_io_slaves_0_w_bits_last;
  assign io_deviceTree_w_bits_data = mmio_ic_io_slaves_0_w_bits_data;
  assign io_deviceTree_w_valid = mmio_ic_io_slaves_0_w_valid;
  assign io_deviceTree_aw_bits_user = mmio_ic_io_slaves_0_aw_bits_user;
  assign io_deviceTree_aw_bits_id = mmio_ic_io_slaves_0_aw_bits_id;
  assign io_deviceTree_aw_bits_region = mmio_ic_io_slaves_0_aw_bits_region;
  assign io_deviceTree_aw_bits_qos = mmio_ic_io_slaves_0_aw_bits_qos;
  assign io_deviceTree_aw_bits_prot = mmio_ic_io_slaves_0_aw_bits_prot;
  assign io_deviceTree_aw_bits_cache = mmio_ic_io_slaves_0_aw_bits_cache;
  assign io_deviceTree_aw_bits_lock = mmio_ic_io_slaves_0_aw_bits_lock;
  assign io_deviceTree_aw_bits_burst = mmio_ic_io_slaves_0_aw_bits_burst;
  assign io_deviceTree_aw_bits_size = mmio_ic_io_slaves_0_aw_bits_size;
  assign io_deviceTree_aw_bits_len = mmio_ic_io_slaves_0_aw_bits_len;
  assign io_deviceTree_aw_bits_addr = mmio_ic_io_slaves_0_aw_bits_addr;
  assign io_deviceTree_aw_valid = mmio_ic_io_slaves_0_aw_valid;
  assign io_scr_resp_ready = scr_conv_io_smi_resp_ready;
  assign io_scr_req_bits_data = scr_conv_io_smi_req_bits_data;
  assign io_scr_req_bits_addr = scr_conv_io_smi_req_bits_addr;
  assign io_scr_req_bits_rw = scr_conv_io_smi_req_bits_rw;
  assign io_scr_req_valid = scr_conv_io_smi_req_valid;
  assign io_csr_0_resp_ready = SmiIONastiIOConverter_io_smi_resp_ready;
  assign io_csr_0_req_bits_data = SmiIONastiIOConverter_io_smi_req_bits_data;
  assign io_csr_0_req_bits_addr = SmiIONastiIOConverter_io_smi_req_bits_addr;
  assign io_csr_0_req_bits_rw = SmiIONastiIOConverter_io_smi_req_bits_rw;
  assign io_csr_0_req_valid = SmiIONastiIOConverter_io_smi_req_valid;
  assign io_mem_backup_req_valid = 1'h0;
  assign io_mem_0_r_ready = mem_ic_io_slaves_0_r_ready;
  assign io_mem_0_ar_bits_user = mem_ic_io_slaves_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = mem_ic_io_slaves_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = mem_ic_io_slaves_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = mem_ic_io_slaves_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = mem_ic_io_slaves_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = mem_ic_io_slaves_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = mem_ic_io_slaves_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = mem_ic_io_slaves_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = mem_ic_io_slaves_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = mem_ic_io_slaves_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = mem_ic_io_slaves_0_ar_bits_addr;
  assign io_mem_0_ar_valid = mem_ic_io_slaves_0_ar_valid;
  assign io_mem_0_b_ready = mem_ic_io_slaves_0_b_ready;
  assign io_mem_0_w_bits_user = mem_ic_io_slaves_0_w_bits_user;
  assign io_mem_0_w_bits_strb = mem_ic_io_slaves_0_w_bits_strb;
  assign io_mem_0_w_bits_last = mem_ic_io_slaves_0_w_bits_last;
  assign io_mem_0_w_bits_data = mem_ic_io_slaves_0_w_bits_data;
  assign io_mem_0_w_valid = mem_ic_io_slaves_0_w_valid;
  assign io_mem_0_aw_bits_user = mem_ic_io_slaves_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = mem_ic_io_slaves_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = mem_ic_io_slaves_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = mem_ic_io_slaves_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = mem_ic_io_slaves_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = mem_ic_io_slaves_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = mem_ic_io_slaves_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = mem_ic_io_slaves_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = mem_ic_io_slaves_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = mem_ic_io_slaves_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = mem_ic_io_slaves_0_aw_bits_addr;
  assign io_mem_0_aw_valid = mem_ic_io_slaves_0_aw_valid;
  assign io_htif_uncached_grant_bits_data = ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  assign io_htif_uncached_grant_bits_g_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  assign io_htif_uncached_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  assign io_htif_uncached_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  assign io_htif_uncached_grant_bits_client_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  assign io_htif_uncached_grant_bits_addr_beat = ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  assign io_htif_uncached_grant_valid = ClientTileLinkIOWrapper_1_io_in_grant_valid;
  assign io_htif_uncached_acquire_ready = ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  assign io_tiles_uncached_0_grant_bits_data = ClientTileLinkIOWrapper_io_in_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = ClientTileLinkIOWrapper_io_in_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = ClientTileLinkIOWrapper_io_in_acquire_ready;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_0_acquire_ready;
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_in_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_in_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper_1(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_1_io_in_acquire_ready ),
       .io_in_acquire_valid( io_htif_uncached_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_htif_uncached_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_htif_uncached_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_htif_uncached_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_htif_uncached_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_htif_uncached_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_htif_uncached_acquire_bits_union ),
       .io_in_acquire_bits_data( io_htif_uncached_acquire_bits_data ),
       .io_in_grant_ready( io_htif_uncached_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_1_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_1_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  RocketChipTileLinkCrossbar l1tol2net(.clk(clk), .reset(reset),
       .io_clients_2_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_clients_2_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_clients_2_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_clients_2_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_clients_2_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_clients_2_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_clients_2_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_clients_2_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_clients_2_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_clients_2_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_clients_2_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_clients_2_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_clients_2_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_clients_2_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_clients_2_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_clients_2_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_clients_2_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_clients_2_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_clients_2_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_clients_2_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_clients_2_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_clients_2_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_clients_2_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid ),
       //.io_clients_2_release_bits_addr_beat(  )
       //.io_clients_2_release_bits_addr_block(  )
       //.io_clients_2_release_bits_client_xact_id(  )
       //.io_clients_2_release_bits_voluntary(  )
       //.io_clients_2_release_bits_r_type(  )
       //.io_clients_2_release_bits_data(  )
       .io_clients_1_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_clients_1_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_clients_1_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_clients_1_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_clients_1_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_clients_1_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_clients_1_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_clients_1_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_clients_1_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_clients_1_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_clients_1_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_clients_1_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_clients_1_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_clients_1_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_clients_1_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_clients_1_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_clients_1_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_clients_1_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_clients_1_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( ClientTileLinkIOWrapper_io_out_release_valid ),
       //.io_clients_1_release_bits_addr_beat(  )
       //.io_clients_1_release_bits_addr_block(  )
       //.io_clients_1_release_bits_client_xact_id(  )
       //.io_clients_1_release_bits_voluntary(  )
       //.io_clients_1_release_bits_r_type(  )
       //.io_clients_1_release_bits_data(  )
       .io_clients_0_acquire_ready( l1tol2net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_clients_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_clients_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_clients_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_clients_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_clients_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_clients_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_clients_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_clients_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_clients_0_grant_valid( l1tol2net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_addr_beat( l1tol2net_io_clients_0_grant_bits_addr_beat ),
       .io_clients_0_grant_bits_client_xact_id( l1tol2net_io_clients_0_grant_bits_client_xact_id ),
       .io_clients_0_grant_bits_manager_xact_id( l1tol2net_io_clients_0_grant_bits_manager_xact_id ),
       .io_clients_0_grant_bits_is_builtin_type( l1tol2net_io_clients_0_grant_bits_is_builtin_type ),
       .io_clients_0_grant_bits_g_type( l1tol2net_io_clients_0_grant_bits_g_type ),
       .io_clients_0_grant_bits_data( l1tol2net_io_clients_0_grant_bits_data ),
       .io_clients_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_clients_0_probe_valid( l1tol2net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_addr_block( l1tol2net_io_clients_0_probe_bits_addr_block ),
       .io_clients_0_probe_bits_p_type( l1tol2net_io_clients_0_probe_bits_p_type ),
       .io_clients_0_release_ready( l1tol2net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_clients_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_clients_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_clients_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_clients_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_clients_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_clients_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_managers_1_acquire_ready( mmioManager_io_inner_acquire_ready ),
       .io_managers_1_acquire_valid( l1tol2net_io_managers_1_acquire_valid ),
       .io_managers_1_acquire_bits_addr_block( l1tol2net_io_managers_1_acquire_bits_addr_block ),
       .io_managers_1_acquire_bits_client_xact_id( l1tol2net_io_managers_1_acquire_bits_client_xact_id ),
       .io_managers_1_acquire_bits_addr_beat( l1tol2net_io_managers_1_acquire_bits_addr_beat ),
       .io_managers_1_acquire_bits_is_builtin_type( l1tol2net_io_managers_1_acquire_bits_is_builtin_type ),
       .io_managers_1_acquire_bits_a_type( l1tol2net_io_managers_1_acquire_bits_a_type ),
       .io_managers_1_acquire_bits_union( l1tol2net_io_managers_1_acquire_bits_union ),
       .io_managers_1_acquire_bits_data( l1tol2net_io_managers_1_acquire_bits_data ),
       .io_managers_1_acquire_bits_client_id( l1tol2net_io_managers_1_acquire_bits_client_id ),
       .io_managers_1_grant_ready( l1tol2net_io_managers_1_grant_ready ),
       .io_managers_1_grant_valid( mmioManager_io_inner_grant_valid ),
       .io_managers_1_grant_bits_addr_beat( mmioManager_io_inner_grant_bits_addr_beat ),
       .io_managers_1_grant_bits_client_xact_id( mmioManager_io_inner_grant_bits_client_xact_id ),
       .io_managers_1_grant_bits_manager_xact_id( mmioManager_io_inner_grant_bits_manager_xact_id ),
       .io_managers_1_grant_bits_is_builtin_type( mmioManager_io_inner_grant_bits_is_builtin_type ),
       .io_managers_1_grant_bits_g_type( mmioManager_io_inner_grant_bits_g_type ),
       .io_managers_1_grant_bits_data( mmioManager_io_inner_grant_bits_data ),
       .io_managers_1_grant_bits_client_id( mmioManager_io_inner_grant_bits_client_id ),
       .io_managers_1_finish_ready( mmioManager_io_inner_finish_ready ),
       .io_managers_1_finish_valid( l1tol2net_io_managers_1_finish_valid ),
       .io_managers_1_finish_bits_manager_xact_id( l1tol2net_io_managers_1_finish_bits_manager_xact_id ),
       .io_managers_1_probe_ready( l1tol2net_io_managers_1_probe_ready ),
       .io_managers_1_probe_valid( mmioManager_io_inner_probe_valid ),
       //.io_managers_1_probe_bits_addr_block(  )
       //.io_managers_1_probe_bits_p_type(  )
       //.io_managers_1_probe_bits_client_id(  )
       .io_managers_1_release_ready( mmioManager_io_inner_release_ready ),
       .io_managers_1_release_valid( l1tol2net_io_managers_1_release_valid ),
       .io_managers_1_release_bits_addr_beat( l1tol2net_io_managers_1_release_bits_addr_beat ),
       .io_managers_1_release_bits_addr_block( l1tol2net_io_managers_1_release_bits_addr_block ),
       .io_managers_1_release_bits_client_xact_id( l1tol2net_io_managers_1_release_bits_client_xact_id ),
       .io_managers_1_release_bits_voluntary( l1tol2net_io_managers_1_release_bits_voluntary ),
       .io_managers_1_release_bits_r_type( l1tol2net_io_managers_1_release_bits_r_type ),
       .io_managers_1_release_bits_data( l1tol2net_io_managers_1_release_bits_data ),
       .io_managers_1_release_bits_client_id( l1tol2net_io_managers_1_release_bits_client_id ),
       .io_managers_0_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_managers_0_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_managers_0_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_managers_0_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_managers_0_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_managers_0_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_managers_0_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_managers_0_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_managers_0_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_managers_0_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_managers_0_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_managers_0_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_managers_0_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_managers_0_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_managers_0_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_managers_0_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_managers_0_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_managers_0_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_managers_0_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_managers_0_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_managers_0_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_managers_0_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_managers_0_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_managers_0_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_managers_0_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_managers_0_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_managers_0_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_managers_0_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_managers_0_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_managers_0_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_managers_0_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_managers_0_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign l1tol2net.io_clients_2_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_data = {4{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_data = {4{$random}};
    assign l1tol2net.io_managers_1_probe_bits_addr_block = {1{$random}};
    assign l1tol2net.io_managers_1_probe_bits_p_type = {1{$random}};
    assign l1tol2net.io_managers_1_probe_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  L2BroadcastHub L2BroadcastHub(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_inner_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_inner_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_inner_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_inner_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_inner_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_inner_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_inner_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_inner_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_inner_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_inner_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_inner_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_inner_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_inner_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_inner_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_outer_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data )
  );
  MMIOTileLinkManager mmioManager(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( mmioManager_io_inner_acquire_ready ),
       .io_inner_acquire_valid( l1tol2net_io_managers_1_acquire_valid ),
       .io_inner_acquire_bits_addr_block( l1tol2net_io_managers_1_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( l1tol2net_io_managers_1_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( l1tol2net_io_managers_1_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( l1tol2net_io_managers_1_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( l1tol2net_io_managers_1_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( l1tol2net_io_managers_1_acquire_bits_union ),
       .io_inner_acquire_bits_data( l1tol2net_io_managers_1_acquire_bits_data ),
       .io_inner_acquire_bits_client_id( l1tol2net_io_managers_1_acquire_bits_client_id ),
       .io_inner_grant_ready( l1tol2net_io_managers_1_grant_ready ),
       .io_inner_grant_valid( mmioManager_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( mmioManager_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( mmioManager_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( mmioManager_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( mmioManager_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( mmioManager_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( mmioManager_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( mmioManager_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( mmioManager_io_inner_finish_ready ),
       .io_inner_finish_valid( l1tol2net_io_managers_1_finish_valid ),
       .io_inner_finish_bits_manager_xact_id( l1tol2net_io_managers_1_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( l1tol2net_io_managers_1_probe_ready ),
       .io_inner_probe_valid( mmioManager_io_inner_probe_valid ),
       //.io_inner_probe_bits_addr_block(  )
       //.io_inner_probe_bits_p_type(  )
       //.io_inner_probe_bits_client_id(  )
       .io_inner_release_ready( mmioManager_io_inner_release_ready ),
       .io_inner_release_valid( l1tol2net_io_managers_1_release_valid ),
       .io_inner_release_bits_addr_beat( l1tol2net_io_managers_1_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( l1tol2net_io_managers_1_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( l1tol2net_io_managers_1_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( l1tol2net_io_managers_1_release_bits_voluntary ),
       .io_inner_release_bits_r_type( l1tol2net_io_managers_1_release_bits_r_type ),
       .io_inner_release_bits_data( l1tol2net_io_managers_1_release_bits_data ),
       .io_inner_release_bits_client_id( l1tol2net_io_managers_1_release_bits_client_id ),
       //.io_incoherent_0(  )
       .io_outer_acquire_ready( mmio_narrow_io_in_acquire_ready ),
       .io_outer_acquire_valid( mmioManager_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( mmioManager_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( mmioManager_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( mmioManager_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( mmioManager_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( mmioManager_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( mmioManager_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( mmioManager_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( mmioManager_io_outer_grant_ready ),
       .io_outer_grant_valid( mmio_narrow_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( mmio_narrow_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( mmio_narrow_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( mmio_narrow_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( mmio_narrow_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( mmio_narrow_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( mmio_narrow_io_in_grant_bits_data )
  );
  NastiRecursiveInterconnect_1 mmio_ic(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( mmio_ic_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( rtc_io_aw_valid ),
       .io_masters_1_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_masters_1_aw_bits_len( rtc_io_aw_bits_len ),
       .io_masters_1_aw_bits_size( rtc_io_aw_bits_size ),
       .io_masters_1_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_masters_1_aw_bits_region( rtc_io_aw_bits_region ),
       .io_masters_1_aw_bits_id( rtc_io_aw_bits_id ),
       .io_masters_1_aw_bits_user( rtc_io_aw_bits_user ),
       .io_masters_1_w_ready( mmio_ic_io_masters_1_w_ready ),
       .io_masters_1_w_valid( rtc_io_w_valid ),
       .io_masters_1_w_bits_data( rtc_io_w_bits_data ),
       .io_masters_1_w_bits_last( rtc_io_w_bits_last ),
       .io_masters_1_w_bits_strb( rtc_io_w_bits_strb ),
       .io_masters_1_w_bits_user( rtc_io_w_bits_user ),
       .io_masters_1_b_ready( rtc_io_b_ready ),
       .io_masters_1_b_valid( mmio_ic_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( mmio_ic_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( mmio_ic_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( mmio_ic_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( mmio_ic_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( rtc_io_ar_valid ),
       //.io_masters_1_ar_bits_addr(  )
       //.io_masters_1_ar_bits_len(  )
       //.io_masters_1_ar_bits_size(  )
       //.io_masters_1_ar_bits_burst(  )
       //.io_masters_1_ar_bits_lock(  )
       //.io_masters_1_ar_bits_cache(  )
       //.io_masters_1_ar_bits_prot(  )
       //.io_masters_1_ar_bits_qos(  )
       //.io_masters_1_ar_bits_region(  )
       //.io_masters_1_ar_bits_id(  )
       //.io_masters_1_ar_bits_user(  )
       .io_masters_1_r_ready( rtc_io_r_ready ),
       .io_masters_1_r_valid( mmio_ic_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( mmio_ic_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( mmio_ic_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( mmio_ic_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( mmio_ic_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( mmio_ic_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( mmio_ic_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( Queue_6_io_deq_valid ),
       .io_masters_0_aw_bits_addr( Queue_6_io_deq_bits_addr ),
       .io_masters_0_aw_bits_len( Queue_6_io_deq_bits_len ),
       .io_masters_0_aw_bits_size( Queue_6_io_deq_bits_size ),
       .io_masters_0_aw_bits_burst( Queue_6_io_deq_bits_burst ),
       .io_masters_0_aw_bits_lock( Queue_6_io_deq_bits_lock ),
       .io_masters_0_aw_bits_cache( Queue_6_io_deq_bits_cache ),
       .io_masters_0_aw_bits_prot( Queue_6_io_deq_bits_prot ),
       .io_masters_0_aw_bits_qos( Queue_6_io_deq_bits_qos ),
       .io_masters_0_aw_bits_region( Queue_6_io_deq_bits_region ),
       .io_masters_0_aw_bits_id( Queue_6_io_deq_bits_id ),
       .io_masters_0_aw_bits_user( Queue_6_io_deq_bits_user ),
       .io_masters_0_w_ready( mmio_ic_io_masters_0_w_ready ),
       .io_masters_0_w_valid( Queue_7_io_deq_valid ),
       .io_masters_0_w_bits_data( Queue_7_io_deq_bits_data ),
       .io_masters_0_w_bits_last( Queue_7_io_deq_bits_last ),
       .io_masters_0_w_bits_strb( Queue_7_io_deq_bits_strb ),
       .io_masters_0_w_bits_user( Queue_7_io_deq_bits_user ),
       .io_masters_0_b_ready( Queue_9_io_enq_ready ),
       .io_masters_0_b_valid( mmio_ic_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( mmio_ic_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( mmio_ic_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( mmio_ic_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( mmio_ic_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( Queue_5_io_deq_valid ),
       .io_masters_0_ar_bits_addr( Queue_5_io_deq_bits_addr ),
       .io_masters_0_ar_bits_len( Queue_5_io_deq_bits_len ),
       .io_masters_0_ar_bits_size( Queue_5_io_deq_bits_size ),
       .io_masters_0_ar_bits_burst( Queue_5_io_deq_bits_burst ),
       .io_masters_0_ar_bits_lock( Queue_5_io_deq_bits_lock ),
       .io_masters_0_ar_bits_cache( Queue_5_io_deq_bits_cache ),
       .io_masters_0_ar_bits_prot( Queue_5_io_deq_bits_prot ),
       .io_masters_0_ar_bits_qos( Queue_5_io_deq_bits_qos ),
       .io_masters_0_ar_bits_region( Queue_5_io_deq_bits_region ),
       .io_masters_0_ar_bits_id( Queue_5_io_deq_bits_id ),
       .io_masters_0_ar_bits_user( Queue_5_io_deq_bits_user ),
       .io_masters_0_r_ready( Queue_8_io_enq_ready ),
       .io_masters_0_r_valid( mmio_ic_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( mmio_ic_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( mmio_ic_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( mmio_ic_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( mmio_ic_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( mmio_ic_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( scr_conv_io_nasti_aw_ready ),
       .io_slaves_2_aw_valid( mmio_ic_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( mmio_ic_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( mmio_ic_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( mmio_ic_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( mmio_ic_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( mmio_ic_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( mmio_ic_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( mmio_ic_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( mmio_ic_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( mmio_ic_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( mmio_ic_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( mmio_ic_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( scr_conv_io_nasti_w_ready ),
       .io_slaves_2_w_valid( mmio_ic_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( mmio_ic_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( mmio_ic_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( mmio_ic_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( mmio_ic_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( mmio_ic_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( scr_conv_io_nasti_b_valid ),
       .io_slaves_2_b_bits_resp( scr_conv_io_nasti_b_bits_resp ),
       .io_slaves_2_b_bits_id( scr_conv_io_nasti_b_bits_id ),
       .io_slaves_2_b_bits_user( scr_conv_io_nasti_b_bits_user ),
       .io_slaves_2_ar_ready( scr_conv_io_nasti_ar_ready ),
       .io_slaves_2_ar_valid( mmio_ic_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( mmio_ic_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( mmio_ic_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( mmio_ic_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( mmio_ic_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( mmio_ic_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( mmio_ic_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( mmio_ic_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( mmio_ic_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( mmio_ic_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( mmio_ic_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( mmio_ic_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( mmio_ic_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( scr_conv_io_nasti_r_valid ),
       .io_slaves_2_r_bits_resp( scr_conv_io_nasti_r_bits_resp ),
       .io_slaves_2_r_bits_data( scr_conv_io_nasti_r_bits_data ),
       .io_slaves_2_r_bits_last( scr_conv_io_nasti_r_bits_last ),
       .io_slaves_2_r_bits_id( scr_conv_io_nasti_r_bits_id ),
       .io_slaves_2_r_bits_user( scr_conv_io_nasti_r_bits_user ),
       .io_slaves_1_aw_ready( SmiIONastiIOConverter_io_nasti_aw_ready ),
       .io_slaves_1_aw_valid( mmio_ic_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( mmio_ic_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( mmio_ic_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( mmio_ic_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( mmio_ic_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( mmio_ic_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( mmio_ic_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( mmio_ic_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( mmio_ic_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( mmio_ic_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( mmio_ic_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( mmio_ic_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( SmiIONastiIOConverter_io_nasti_w_ready ),
       .io_slaves_1_w_valid( mmio_ic_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( mmio_ic_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( mmio_ic_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( mmio_ic_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( mmio_ic_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( mmio_ic_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( SmiIONastiIOConverter_io_nasti_b_valid ),
       .io_slaves_1_b_bits_resp( SmiIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_slaves_1_b_bits_id( SmiIONastiIOConverter_io_nasti_b_bits_id ),
       .io_slaves_1_b_bits_user( SmiIONastiIOConverter_io_nasti_b_bits_user ),
       .io_slaves_1_ar_ready( SmiIONastiIOConverter_io_nasti_ar_ready ),
       .io_slaves_1_ar_valid( mmio_ic_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( mmio_ic_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( mmio_ic_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( mmio_ic_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( mmio_ic_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( mmio_ic_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( mmio_ic_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( mmio_ic_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( mmio_ic_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( mmio_ic_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( mmio_ic_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( mmio_ic_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( mmio_ic_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( SmiIONastiIOConverter_io_nasti_r_valid ),
       .io_slaves_1_r_bits_resp( SmiIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_slaves_1_r_bits_data( SmiIONastiIOConverter_io_nasti_r_bits_data ),
       .io_slaves_1_r_bits_last( SmiIONastiIOConverter_io_nasti_r_bits_last ),
       .io_slaves_1_r_bits_id( SmiIONastiIOConverter_io_nasti_r_bits_id ),
       .io_slaves_1_r_bits_user( SmiIONastiIOConverter_io_nasti_r_bits_user ),
       .io_slaves_0_aw_ready( io_deviceTree_aw_ready ),
       .io_slaves_0_aw_valid( mmio_ic_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( mmio_ic_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( mmio_ic_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( mmio_ic_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( mmio_ic_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( mmio_ic_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( mmio_ic_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( mmio_ic_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( mmio_ic_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( mmio_ic_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( mmio_ic_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( mmio_ic_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_deviceTree_w_ready ),
       .io_slaves_0_w_valid( mmio_ic_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( mmio_ic_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( mmio_ic_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( mmio_ic_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( mmio_ic_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( mmio_ic_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_deviceTree_b_valid ),
       .io_slaves_0_b_bits_resp( io_deviceTree_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_deviceTree_b_bits_id ),
       .io_slaves_0_b_bits_user( io_deviceTree_b_bits_user ),
       .io_slaves_0_ar_ready( io_deviceTree_ar_ready ),
       .io_slaves_0_ar_valid( mmio_ic_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( mmio_ic_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( mmio_ic_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( mmio_ic_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( mmio_ic_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( mmio_ic_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( mmio_ic_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( mmio_ic_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( mmio_ic_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( mmio_ic_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( mmio_ic_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( mmio_ic_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( mmio_ic_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_deviceTree_r_valid ),
       .io_slaves_0_r_bits_resp( io_deviceTree_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_deviceTree_r_bits_data ),
       .io_slaves_0_r_bits_last( io_deviceTree_r_bits_last ),
       .io_slaves_0_r_bits_id( io_deviceTree_r_bits_id ),
       .io_slaves_0_r_bits_user( io_deviceTree_r_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign mmio_ic.io_masters_1_ar_bits_addr = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_len = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_size = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_burst = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_lock = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_cache = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_prot = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_qos = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_region = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_id = {1{$random}};
    assign mmio_ic.io_masters_1_ar_bits_user = {1{$random}};
// synthesis translate_on
`endif
  NastiMemoryInterconnect mem_ic(
       .io_masters_0_aw_ready( mem_ic_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( Queue_1_io_deq_valid ),
       .io_masters_0_aw_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_masters_0_aw_bits_len( Queue_1_io_deq_bits_len ),
       .io_masters_0_aw_bits_size( Queue_1_io_deq_bits_size ),
       .io_masters_0_aw_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_masters_0_aw_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_masters_0_aw_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_masters_0_aw_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_masters_0_aw_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_masters_0_aw_bits_region( Queue_1_io_deq_bits_region ),
       .io_masters_0_aw_bits_id( Queue_1_io_deq_bits_id ),
       .io_masters_0_aw_bits_user( Queue_1_io_deq_bits_user ),
       .io_masters_0_w_ready( mem_ic_io_masters_0_w_ready ),
       .io_masters_0_w_valid( Queue_2_io_deq_valid ),
       .io_masters_0_w_bits_data( Queue_2_io_deq_bits_data ),
       .io_masters_0_w_bits_last( Queue_2_io_deq_bits_last ),
       .io_masters_0_w_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_masters_0_w_bits_user( Queue_2_io_deq_bits_user ),
       .io_masters_0_b_ready( Queue_4_io_enq_ready ),
       .io_masters_0_b_valid( mem_ic_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( mem_ic_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( mem_ic_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( mem_ic_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( mem_ic_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( Queue_io_deq_valid ),
       .io_masters_0_ar_bits_addr( Queue_io_deq_bits_addr ),
       .io_masters_0_ar_bits_len( Queue_io_deq_bits_len ),
       .io_masters_0_ar_bits_size( Queue_io_deq_bits_size ),
       .io_masters_0_ar_bits_burst( Queue_io_deq_bits_burst ),
       .io_masters_0_ar_bits_lock( Queue_io_deq_bits_lock ),
       .io_masters_0_ar_bits_cache( Queue_io_deq_bits_cache ),
       .io_masters_0_ar_bits_prot( Queue_io_deq_bits_prot ),
       .io_masters_0_ar_bits_qos( Queue_io_deq_bits_qos ),
       .io_masters_0_ar_bits_region( Queue_io_deq_bits_region ),
       .io_masters_0_ar_bits_id( Queue_io_deq_bits_id ),
       .io_masters_0_ar_bits_user( Queue_io_deq_bits_user ),
       .io_masters_0_r_ready( Queue_3_io_enq_ready ),
       .io_masters_0_r_valid( mem_ic_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( mem_ic_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( mem_ic_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( mem_ic_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( mem_ic_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( mem_ic_io_masters_0_r_bits_user ),
       .io_slaves_0_aw_ready( io_mem_0_aw_ready ),
       .io_slaves_0_aw_valid( mem_ic_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( mem_ic_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( mem_ic_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( mem_ic_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( mem_ic_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( mem_ic_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( mem_ic_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( mem_ic_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( mem_ic_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( mem_ic_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( mem_ic_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( mem_ic_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_mem_0_w_ready ),
       .io_slaves_0_w_valid( mem_ic_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( mem_ic_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( mem_ic_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( mem_ic_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( mem_ic_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( mem_ic_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_mem_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_mem_0_ar_ready ),
       .io_slaves_0_ar_valid( mem_ic_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( mem_ic_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( mem_ic_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( mem_ic_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( mem_ic_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( mem_ic_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( mem_ic_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( mem_ic_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( mem_ic_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( mem_ic_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( mem_ic_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( mem_ic_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( mem_ic_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_mem_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_mem_0_r_bits_user )
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper(.clk(clk), .reset(reset),
       .io_in_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkEnqueuer_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkEnqueuer_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkEnqueuer_io_outer_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkEnqueuer_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_in_probe_ready( ClientTileLinkEnqueuer_io_outer_probe_ready ),
       .io_in_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_in_probe_bits_addr_block(  )
       //.io_in_probe_bits_p_type(  )
       .io_in_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_in_release_valid( ClientTileLinkEnqueuer_io_outer_release_valid ),
       .io_in_release_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat ),
       .io_in_release_bits_addr_block( ClientTileLinkEnqueuer_io_outer_release_bits_addr_block ),
       .io_in_release_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id ),
       .io_in_release_bits_voluntary( ClientTileLinkEnqueuer_io_outer_release_bits_voluntary ),
       .io_in_release_bits_r_type( ClientTileLinkEnqueuer_io_outer_release_bits_r_type ),
       .io_in_release_bits_data( ClientTileLinkEnqueuer_io_outer_release_bits_data ),
       .io_out_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_out_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_out_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_out_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data )
  );
  TileLinkIONarrower TileLinkIONarrower(.clk(clk), .reset(reset),
       .io_in_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_in_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data ),
       .io_out_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_out_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_out_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_out_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_out_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_out_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data )
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_tl_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_tl_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_tl_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_tl_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_tl_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data ),
       .io_nasti_aw_ready( Queue_1_io_enq_ready ),
       .io_nasti_aw_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_nasti_aw_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_nasti_aw_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_nasti_aw_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_nasti_aw_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_nasti_aw_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_nasti_aw_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_nasti_aw_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_nasti_aw_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_nasti_aw_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_nasti_aw_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_nasti_aw_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_nasti_w_ready( Queue_2_io_enq_ready ),
       .io_nasti_w_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_nasti_w_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_nasti_w_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_nasti_w_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_nasti_w_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_nasti_b_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_nasti_b_valid( Queue_4_io_deq_valid ),
       .io_nasti_b_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_nasti_b_bits_id( Queue_4_io_deq_bits_id ),
       .io_nasti_b_bits_user( Queue_4_io_deq_bits_user ),
       .io_nasti_ar_ready( Queue_io_enq_ready ),
       .io_nasti_ar_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_nasti_ar_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_nasti_ar_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_nasti_ar_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_nasti_ar_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_nasti_ar_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_nasti_ar_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_nasti_ar_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_nasti_ar_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_nasti_ar_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_nasti_ar_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_nasti_ar_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_nasti_r_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_nasti_r_valid( Queue_3_io_deq_valid ),
       .io_nasti_r_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_nasti_r_bits_data( Queue_3_io_deq_bits_data ),
       .io_nasti_r_bits_last( Queue_3_io_deq_bits_last ),
       .io_nasti_r_bits_id( Queue_3_io_deq_bits_id ),
       .io_nasti_r_bits_user( Queue_3_io_deq_bits_user )
  );
  ClientTileLinkIOWrapper_1 ClientTileLinkIOWrapper_2(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_in_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_in_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data ),
       .io_out_acquire_ready( ClientTileLinkEnqueuer_io_inner_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_out_grant_valid( ClientTileLinkEnqueuer_io_inner_grant_valid ),
       .io_out_grant_bits_addr_beat( ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( ClientTileLinkEnqueuer_io_inner_grant_bits_g_type ),
       .io_out_grant_bits_data( ClientTileLinkEnqueuer_io_inner_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_out_probe_valid( ClientTileLinkEnqueuer_io_inner_probe_valid ),
       .io_out_probe_bits_addr_block( ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( ClientTileLinkEnqueuer_io_inner_probe_bits_p_type ),
       .io_out_release_ready( ClientTileLinkEnqueuer_io_inner_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer(
       .io_inner_acquire_ready( ClientTileLinkEnqueuer_io_inner_acquire_ready ),
       .io_inner_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_inner_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_inner_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_inner_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_inner_grant_valid( ClientTileLinkEnqueuer_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( ClientTileLinkEnqueuer_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( ClientTileLinkEnqueuer_io_inner_grant_bits_data ),
       .io_inner_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_inner_probe_valid( ClientTileLinkEnqueuer_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( ClientTileLinkEnqueuer_io_inner_probe_bits_p_type ),
       .io_inner_release_ready( ClientTileLinkEnqueuer_io_inner_release_ready ),
       .io_inner_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid ),
       //.io_inner_release_bits_addr_beat(  )
       //.io_inner_release_bits_addr_block(  )
       //.io_inner_release_bits_client_xact_id(  )
       //.io_inner_release_bits_voluntary(  )
       //.io_inner_release_bits_r_type(  )
       //.io_inner_release_bits_data(  )
       .io_outer_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_outer_acquire_valid( ClientTileLinkEnqueuer_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( ClientTileLinkEnqueuer_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( ClientTileLinkEnqueuer_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( ClientTileLinkEnqueuer_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_outer_probe_ready( ClientTileLinkEnqueuer_io_outer_probe_ready ),
       .io_outer_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_outer_probe_bits_addr_block(  )
       //.io_outer_probe_bits_p_type(  )
       .io_outer_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_outer_release_valid( ClientTileLinkEnqueuer_io_outer_release_valid ),
       .io_outer_release_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat ),
       .io_outer_release_bits_addr_block( ClientTileLinkEnqueuer_io_outer_release_bits_addr_block ),
       .io_outer_release_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id ),
       .io_outer_release_bits_voluntary( ClientTileLinkEnqueuer_io_outer_release_bits_voluntary ),
       .io_outer_release_bits_r_type( ClientTileLinkEnqueuer_io_outer_release_bits_r_type ),
       .io_outer_release_bits_data( ClientTileLinkEnqueuer_io_outer_release_bits_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ClientTileLinkEnqueuer.io_inner_release_bits_addr_beat = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_addr_block = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_voluntary = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_r_type = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_data = {4{$random}};
    assign ClientTileLinkEnqueuer.io_outer_probe_bits_addr_block = {1{$random}};
    assign ClientTileLinkEnqueuer.io_outer_probe_bits_p_type = {1{$random}};
// synthesis translate_on
`endif
  Queue_2 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_deq_ready( mem_ic_io_masters_0_ar_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_io_deq_bits_len ),
       .io_deq_bits_size( Queue_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_io_deq_bits_region ),
       .io_deq_bits_id( Queue_io_deq_bits_id ),
       .io_deq_bits_user( Queue_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_2 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_deq_ready( mem_ic_io_masters_0_aw_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_1_io_deq_bits_len ),
       .io_deq_bits_size( Queue_1_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_1_io_deq_bits_region ),
       .io_deq_bits_id( Queue_1_io_deq_bits_id ),
       .io_deq_bits_user( Queue_1_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_enq_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_enq_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_enq_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_deq_ready( mem_ic_io_masters_0_w_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_data( Queue_2_io_deq_bits_data ),
       .io_deq_bits_last( Queue_2_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_2_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( mem_ic_io_masters_0_r_valid ),
       .io_enq_bits_resp( mem_ic_io_masters_0_r_bits_resp ),
       .io_enq_bits_data( mem_ic_io_masters_0_r_bits_data ),
       .io_enq_bits_last( mem_ic_io_masters_0_r_bits_last ),
       .io_enq_bits_id( mem_ic_io_masters_0_r_bits_id ),
       .io_enq_bits_user( mem_ic_io_masters_0_r_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_3_io_deq_bits_data ),
       .io_deq_bits_last( Queue_3_io_deq_bits_last ),
       .io_deq_bits_id( Queue_3_io_deq_bits_id ),
       .io_deq_bits_user( Queue_3_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( mem_ic_io_masters_0_b_valid ),
       .io_enq_bits_resp( mem_ic_io_masters_0_b_bits_resp ),
       .io_enq_bits_id( mem_ic_io_masters_0_b_bits_id ),
       .io_enq_bits_user( mem_ic_io_masters_0_b_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_4_io_deq_bits_id ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  TileLinkIONarrower mmio_narrow(.clk(clk), .reset(reset),
       .io_in_acquire_ready( mmio_narrow_io_in_acquire_ready ),
       .io_in_acquire_valid( mmioManager_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( mmioManager_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( mmioManager_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( mmioManager_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( mmioManager_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( mmioManager_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( mmioManager_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( mmioManager_io_outer_acquire_bits_data ),
       .io_in_grant_ready( mmioManager_io_outer_grant_ready ),
       .io_in_grant_valid( mmio_narrow_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( mmio_narrow_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( mmio_narrow_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( mmio_narrow_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( mmio_narrow_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( mmio_narrow_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( mmio_narrow_io_in_grant_bits_data ),
       .io_out_acquire_ready( mmio_conv_io_tl_acquire_ready ),
       .io_out_acquire_valid( mmio_narrow_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( mmio_narrow_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( mmio_narrow_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( mmio_narrow_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( mmio_narrow_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( mmio_narrow_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( mmio_narrow_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( mmio_narrow_io_out_acquire_bits_data ),
       .io_out_grant_ready( mmio_narrow_io_out_grant_ready ),
       .io_out_grant_valid( mmio_conv_io_tl_grant_valid ),
       .io_out_grant_bits_addr_beat( mmio_conv_io_tl_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( mmio_conv_io_tl_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( mmio_conv_io_tl_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( mmio_conv_io_tl_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( mmio_conv_io_tl_grant_bits_g_type ),
       .io_out_grant_bits_data( mmio_conv_io_tl_grant_bits_data )
  );
  NastiIOTileLinkIOConverter mmio_conv(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( mmio_conv_io_tl_acquire_ready ),
       .io_tl_acquire_valid( mmio_narrow_io_out_acquire_valid ),
       .io_tl_acquire_bits_addr_block( mmio_narrow_io_out_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( mmio_narrow_io_out_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( mmio_narrow_io_out_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_is_builtin_type( mmio_narrow_io_out_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( mmio_narrow_io_out_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( mmio_narrow_io_out_acquire_bits_union ),
       .io_tl_acquire_bits_data( mmio_narrow_io_out_acquire_bits_data ),
       .io_tl_grant_ready( mmio_narrow_io_out_grant_ready ),
       .io_tl_grant_valid( mmio_conv_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( mmio_conv_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_client_xact_id( mmio_conv_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( mmio_conv_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( mmio_conv_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( mmio_conv_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_data( mmio_conv_io_tl_grant_bits_data ),
       .io_nasti_aw_ready( Queue_6_io_enq_ready ),
       .io_nasti_aw_valid( mmio_conv_io_nasti_aw_valid ),
       .io_nasti_aw_bits_addr( mmio_conv_io_nasti_aw_bits_addr ),
       .io_nasti_aw_bits_len( mmio_conv_io_nasti_aw_bits_len ),
       .io_nasti_aw_bits_size( mmio_conv_io_nasti_aw_bits_size ),
       .io_nasti_aw_bits_burst( mmio_conv_io_nasti_aw_bits_burst ),
       .io_nasti_aw_bits_lock( mmio_conv_io_nasti_aw_bits_lock ),
       .io_nasti_aw_bits_cache( mmio_conv_io_nasti_aw_bits_cache ),
       .io_nasti_aw_bits_prot( mmio_conv_io_nasti_aw_bits_prot ),
       .io_nasti_aw_bits_qos( mmio_conv_io_nasti_aw_bits_qos ),
       .io_nasti_aw_bits_region( mmio_conv_io_nasti_aw_bits_region ),
       .io_nasti_aw_bits_id( mmio_conv_io_nasti_aw_bits_id ),
       .io_nasti_aw_bits_user( mmio_conv_io_nasti_aw_bits_user ),
       .io_nasti_w_ready( Queue_7_io_enq_ready ),
       .io_nasti_w_valid( mmio_conv_io_nasti_w_valid ),
       .io_nasti_w_bits_data( mmio_conv_io_nasti_w_bits_data ),
       .io_nasti_w_bits_last( mmio_conv_io_nasti_w_bits_last ),
       .io_nasti_w_bits_strb( mmio_conv_io_nasti_w_bits_strb ),
       .io_nasti_w_bits_user( mmio_conv_io_nasti_w_bits_user ),
       .io_nasti_b_ready( mmio_conv_io_nasti_b_ready ),
       .io_nasti_b_valid( Queue_9_io_deq_valid ),
       .io_nasti_b_bits_resp( Queue_9_io_deq_bits_resp ),
       .io_nasti_b_bits_id( Queue_9_io_deq_bits_id ),
       .io_nasti_b_bits_user( Queue_9_io_deq_bits_user ),
       .io_nasti_ar_ready( Queue_5_io_enq_ready ),
       .io_nasti_ar_valid( mmio_conv_io_nasti_ar_valid ),
       .io_nasti_ar_bits_addr( mmio_conv_io_nasti_ar_bits_addr ),
       .io_nasti_ar_bits_len( mmio_conv_io_nasti_ar_bits_len ),
       .io_nasti_ar_bits_size( mmio_conv_io_nasti_ar_bits_size ),
       .io_nasti_ar_bits_burst( mmio_conv_io_nasti_ar_bits_burst ),
       .io_nasti_ar_bits_lock( mmio_conv_io_nasti_ar_bits_lock ),
       .io_nasti_ar_bits_cache( mmio_conv_io_nasti_ar_bits_cache ),
       .io_nasti_ar_bits_prot( mmio_conv_io_nasti_ar_bits_prot ),
       .io_nasti_ar_bits_qos( mmio_conv_io_nasti_ar_bits_qos ),
       .io_nasti_ar_bits_region( mmio_conv_io_nasti_ar_bits_region ),
       .io_nasti_ar_bits_id( mmio_conv_io_nasti_ar_bits_id ),
       .io_nasti_ar_bits_user( mmio_conv_io_nasti_ar_bits_user ),
       .io_nasti_r_ready( mmio_conv_io_nasti_r_ready ),
       .io_nasti_r_valid( Queue_8_io_deq_valid ),
       .io_nasti_r_bits_resp( Queue_8_io_deq_bits_resp ),
       .io_nasti_r_bits_data( Queue_8_io_deq_bits_data ),
       .io_nasti_r_bits_last( Queue_8_io_deq_bits_last ),
       .io_nasti_r_bits_id( Queue_8_io_deq_bits_id ),
       .io_nasti_r_bits_user( Queue_8_io_deq_bits_user )
  );
  Queue_2 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( mmio_conv_io_nasti_ar_valid ),
       .io_enq_bits_addr( mmio_conv_io_nasti_ar_bits_addr ),
       .io_enq_bits_len( mmio_conv_io_nasti_ar_bits_len ),
       .io_enq_bits_size( mmio_conv_io_nasti_ar_bits_size ),
       .io_enq_bits_burst( mmio_conv_io_nasti_ar_bits_burst ),
       .io_enq_bits_lock( mmio_conv_io_nasti_ar_bits_lock ),
       .io_enq_bits_cache( mmio_conv_io_nasti_ar_bits_cache ),
       .io_enq_bits_prot( mmio_conv_io_nasti_ar_bits_prot ),
       .io_enq_bits_qos( mmio_conv_io_nasti_ar_bits_qos ),
       .io_enq_bits_region( mmio_conv_io_nasti_ar_bits_region ),
       .io_enq_bits_id( mmio_conv_io_nasti_ar_bits_id ),
       .io_enq_bits_user( mmio_conv_io_nasti_ar_bits_user ),
       .io_deq_ready( mmio_ic_io_masters_0_ar_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_addr( Queue_5_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_5_io_deq_bits_len ),
       .io_deq_bits_size( Queue_5_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_5_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_5_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_5_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_5_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_5_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_5_io_deq_bits_region ),
       .io_deq_bits_id( Queue_5_io_deq_bits_id ),
       .io_deq_bits_user( Queue_5_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_2 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( mmio_conv_io_nasti_aw_valid ),
       .io_enq_bits_addr( mmio_conv_io_nasti_aw_bits_addr ),
       .io_enq_bits_len( mmio_conv_io_nasti_aw_bits_len ),
       .io_enq_bits_size( mmio_conv_io_nasti_aw_bits_size ),
       .io_enq_bits_burst( mmio_conv_io_nasti_aw_bits_burst ),
       .io_enq_bits_lock( mmio_conv_io_nasti_aw_bits_lock ),
       .io_enq_bits_cache( mmio_conv_io_nasti_aw_bits_cache ),
       .io_enq_bits_prot( mmio_conv_io_nasti_aw_bits_prot ),
       .io_enq_bits_qos( mmio_conv_io_nasti_aw_bits_qos ),
       .io_enq_bits_region( mmio_conv_io_nasti_aw_bits_region ),
       .io_enq_bits_id( mmio_conv_io_nasti_aw_bits_id ),
       .io_enq_bits_user( mmio_conv_io_nasti_aw_bits_user ),
       .io_deq_ready( mmio_ic_io_masters_0_aw_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_addr( Queue_6_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_6_io_deq_bits_len ),
       .io_deq_bits_size( Queue_6_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_6_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_6_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_6_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_6_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_6_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_6_io_deq_bits_region ),
       .io_deq_bits_id( Queue_6_io_deq_bits_id ),
       .io_deq_bits_user( Queue_6_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( mmio_conv_io_nasti_w_valid ),
       .io_enq_bits_data( mmio_conv_io_nasti_w_bits_data ),
       .io_enq_bits_last( mmio_conv_io_nasti_w_bits_last ),
       .io_enq_bits_strb( mmio_conv_io_nasti_w_bits_strb ),
       .io_enq_bits_user( mmio_conv_io_nasti_w_bits_user ),
       .io_deq_ready( mmio_ic_io_masters_0_w_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_data( Queue_7_io_deq_bits_data ),
       .io_deq_bits_last( Queue_7_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_7_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_7_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( mmio_ic_io_masters_0_r_valid ),
       .io_enq_bits_resp( mmio_ic_io_masters_0_r_bits_resp ),
       .io_enq_bits_data( mmio_ic_io_masters_0_r_bits_data ),
       .io_enq_bits_last( mmio_ic_io_masters_0_r_bits_last ),
       .io_enq_bits_id( mmio_ic_io_masters_0_r_bits_id ),
       .io_enq_bits_user( mmio_ic_io_masters_0_r_bits_user ),
       .io_deq_ready( mmio_conv_io_nasti_r_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_resp( Queue_8_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_8_io_deq_bits_data ),
       .io_deq_bits_last( Queue_8_io_deq_bits_last ),
       .io_deq_bits_id( Queue_8_io_deq_bits_id ),
       .io_deq_bits_user( Queue_8_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( mmio_ic_io_masters_0_b_valid ),
       .io_enq_bits_resp( mmio_ic_io_masters_0_b_bits_resp ),
       .io_enq_bits_id( mmio_ic_io_masters_0_b_bits_id ),
       .io_enq_bits_user( mmio_ic_io_masters_0_b_bits_user ),
       .io_deq_ready( mmio_conv_io_nasti_b_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_resp( Queue_9_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_9_io_deq_bits_id ),
       .io_deq_bits_user( Queue_9_io_deq_bits_user )
       //.io_count(  )
  );
  RTC rtc(.clk(clk), .reset(reset),
       .io_aw_ready( mmio_ic_io_masters_1_aw_ready ),
       .io_aw_valid( rtc_io_aw_valid ),
       .io_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_aw_bits_len( rtc_io_aw_bits_len ),
       .io_aw_bits_size( rtc_io_aw_bits_size ),
       .io_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_aw_bits_region( rtc_io_aw_bits_region ),
       .io_aw_bits_id( rtc_io_aw_bits_id ),
       .io_aw_bits_user( rtc_io_aw_bits_user ),
       .io_w_ready( mmio_ic_io_masters_1_w_ready ),
       .io_w_valid( rtc_io_w_valid ),
       .io_w_bits_data( rtc_io_w_bits_data ),
       .io_w_bits_last( rtc_io_w_bits_last ),
       .io_w_bits_strb( rtc_io_w_bits_strb ),
       .io_w_bits_user( rtc_io_w_bits_user ),
       .io_b_ready( rtc_io_b_ready ),
       .io_b_valid( mmio_ic_io_masters_1_b_valid ),
       .io_b_bits_resp( mmio_ic_io_masters_1_b_bits_resp ),
       .io_b_bits_id( mmio_ic_io_masters_1_b_bits_id ),
       .io_b_bits_user( mmio_ic_io_masters_1_b_bits_user ),
       .io_ar_ready( mmio_ic_io_masters_1_ar_ready ),
       .io_ar_valid( rtc_io_ar_valid ),
       //.io_ar_bits_addr(  )
       //.io_ar_bits_len(  )
       //.io_ar_bits_size(  )
       //.io_ar_bits_burst(  )
       //.io_ar_bits_lock(  )
       //.io_ar_bits_cache(  )
       //.io_ar_bits_prot(  )
       //.io_ar_bits_qos(  )
       //.io_ar_bits_region(  )
       //.io_ar_bits_id(  )
       //.io_ar_bits_user(  )
       .io_r_ready( rtc_io_r_ready ),
       .io_r_valid( mmio_ic_io_masters_1_r_valid ),
       .io_r_bits_resp( mmio_ic_io_masters_1_r_bits_resp ),
       .io_r_bits_data( mmio_ic_io_masters_1_r_bits_data ),
       .io_r_bits_last( mmio_ic_io_masters_1_r_bits_last ),
       .io_r_bits_id( mmio_ic_io_masters_1_r_bits_id ),
       .io_r_bits_user( mmio_ic_io_masters_1_r_bits_user )
  );
  SmiIONastiIOConverter_0 SmiIONastiIOConverter(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( SmiIONastiIOConverter_io_nasti_aw_ready ),
       .io_nasti_aw_valid( mmio_ic_io_slaves_1_aw_valid ),
       .io_nasti_aw_bits_addr( mmio_ic_io_slaves_1_aw_bits_addr ),
       .io_nasti_aw_bits_len( mmio_ic_io_slaves_1_aw_bits_len ),
       .io_nasti_aw_bits_size( mmio_ic_io_slaves_1_aw_bits_size ),
       .io_nasti_aw_bits_burst( mmio_ic_io_slaves_1_aw_bits_burst ),
       .io_nasti_aw_bits_lock( mmio_ic_io_slaves_1_aw_bits_lock ),
       .io_nasti_aw_bits_cache( mmio_ic_io_slaves_1_aw_bits_cache ),
       .io_nasti_aw_bits_prot( mmio_ic_io_slaves_1_aw_bits_prot ),
       .io_nasti_aw_bits_qos( mmio_ic_io_slaves_1_aw_bits_qos ),
       .io_nasti_aw_bits_region( mmio_ic_io_slaves_1_aw_bits_region ),
       .io_nasti_aw_bits_id( mmio_ic_io_slaves_1_aw_bits_id ),
       .io_nasti_aw_bits_user( mmio_ic_io_slaves_1_aw_bits_user ),
       .io_nasti_w_ready( SmiIONastiIOConverter_io_nasti_w_ready ),
       .io_nasti_w_valid( mmio_ic_io_slaves_1_w_valid ),
       .io_nasti_w_bits_data( mmio_ic_io_slaves_1_w_bits_data ),
       .io_nasti_w_bits_last( mmio_ic_io_slaves_1_w_bits_last ),
       .io_nasti_w_bits_strb( mmio_ic_io_slaves_1_w_bits_strb ),
       .io_nasti_w_bits_user( mmio_ic_io_slaves_1_w_bits_user ),
       .io_nasti_b_ready( mmio_ic_io_slaves_1_b_ready ),
       .io_nasti_b_valid( SmiIONastiIOConverter_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( SmiIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( SmiIONastiIOConverter_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( SmiIONastiIOConverter_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( SmiIONastiIOConverter_io_nasti_ar_ready ),
       .io_nasti_ar_valid( mmio_ic_io_slaves_1_ar_valid ),
       .io_nasti_ar_bits_addr( mmio_ic_io_slaves_1_ar_bits_addr ),
       .io_nasti_ar_bits_len( mmio_ic_io_slaves_1_ar_bits_len ),
       .io_nasti_ar_bits_size( mmio_ic_io_slaves_1_ar_bits_size ),
       .io_nasti_ar_bits_burst( mmio_ic_io_slaves_1_ar_bits_burst ),
       .io_nasti_ar_bits_lock( mmio_ic_io_slaves_1_ar_bits_lock ),
       .io_nasti_ar_bits_cache( mmio_ic_io_slaves_1_ar_bits_cache ),
       .io_nasti_ar_bits_prot( mmio_ic_io_slaves_1_ar_bits_prot ),
       .io_nasti_ar_bits_qos( mmio_ic_io_slaves_1_ar_bits_qos ),
       .io_nasti_ar_bits_region( mmio_ic_io_slaves_1_ar_bits_region ),
       .io_nasti_ar_bits_id( mmio_ic_io_slaves_1_ar_bits_id ),
       .io_nasti_ar_bits_user( mmio_ic_io_slaves_1_ar_bits_user ),
       .io_nasti_r_ready( mmio_ic_io_slaves_1_r_ready ),
       .io_nasti_r_valid( SmiIONastiIOConverter_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( SmiIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( SmiIONastiIOConverter_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( SmiIONastiIOConverter_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( SmiIONastiIOConverter_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( SmiIONastiIOConverter_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_csr_0_req_ready ),
       .io_smi_req_valid( SmiIONastiIOConverter_io_smi_req_valid ),
       .io_smi_req_bits_rw( SmiIONastiIOConverter_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( SmiIONastiIOConverter_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( SmiIONastiIOConverter_io_smi_req_bits_data ),
       .io_smi_resp_ready( SmiIONastiIOConverter_io_smi_resp_ready ),
       .io_smi_resp_valid( io_csr_0_resp_valid ),
       .io_smi_resp_bits( io_csr_0_resp_bits )
  );
  SmiIONastiIOConverter_1 scr_conv(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( scr_conv_io_nasti_aw_ready ),
       .io_nasti_aw_valid( mmio_ic_io_slaves_2_aw_valid ),
       .io_nasti_aw_bits_addr( mmio_ic_io_slaves_2_aw_bits_addr ),
       .io_nasti_aw_bits_len( mmio_ic_io_slaves_2_aw_bits_len ),
       .io_nasti_aw_bits_size( mmio_ic_io_slaves_2_aw_bits_size ),
       .io_nasti_aw_bits_burst( mmio_ic_io_slaves_2_aw_bits_burst ),
       .io_nasti_aw_bits_lock( mmio_ic_io_slaves_2_aw_bits_lock ),
       .io_nasti_aw_bits_cache( mmio_ic_io_slaves_2_aw_bits_cache ),
       .io_nasti_aw_bits_prot( mmio_ic_io_slaves_2_aw_bits_prot ),
       .io_nasti_aw_bits_qos( mmio_ic_io_slaves_2_aw_bits_qos ),
       .io_nasti_aw_bits_region( mmio_ic_io_slaves_2_aw_bits_region ),
       .io_nasti_aw_bits_id( mmio_ic_io_slaves_2_aw_bits_id ),
       .io_nasti_aw_bits_user( mmio_ic_io_slaves_2_aw_bits_user ),
       .io_nasti_w_ready( scr_conv_io_nasti_w_ready ),
       .io_nasti_w_valid( mmio_ic_io_slaves_2_w_valid ),
       .io_nasti_w_bits_data( mmio_ic_io_slaves_2_w_bits_data ),
       .io_nasti_w_bits_last( mmio_ic_io_slaves_2_w_bits_last ),
       .io_nasti_w_bits_strb( mmio_ic_io_slaves_2_w_bits_strb ),
       .io_nasti_w_bits_user( mmio_ic_io_slaves_2_w_bits_user ),
       .io_nasti_b_ready( mmio_ic_io_slaves_2_b_ready ),
       .io_nasti_b_valid( scr_conv_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( scr_conv_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( scr_conv_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( scr_conv_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( scr_conv_io_nasti_ar_ready ),
       .io_nasti_ar_valid( mmio_ic_io_slaves_2_ar_valid ),
       .io_nasti_ar_bits_addr( mmio_ic_io_slaves_2_ar_bits_addr ),
       .io_nasti_ar_bits_len( mmio_ic_io_slaves_2_ar_bits_len ),
       .io_nasti_ar_bits_size( mmio_ic_io_slaves_2_ar_bits_size ),
       .io_nasti_ar_bits_burst( mmio_ic_io_slaves_2_ar_bits_burst ),
       .io_nasti_ar_bits_lock( mmio_ic_io_slaves_2_ar_bits_lock ),
       .io_nasti_ar_bits_cache( mmio_ic_io_slaves_2_ar_bits_cache ),
       .io_nasti_ar_bits_prot( mmio_ic_io_slaves_2_ar_bits_prot ),
       .io_nasti_ar_bits_qos( mmio_ic_io_slaves_2_ar_bits_qos ),
       .io_nasti_ar_bits_region( mmio_ic_io_slaves_2_ar_bits_region ),
       .io_nasti_ar_bits_id( mmio_ic_io_slaves_2_ar_bits_id ),
       .io_nasti_ar_bits_user( mmio_ic_io_slaves_2_ar_bits_user ),
       .io_nasti_r_ready( mmio_ic_io_slaves_2_r_ready ),
       .io_nasti_r_valid( scr_conv_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( scr_conv_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( scr_conv_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( scr_conv_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( scr_conv_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( scr_conv_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_scr_req_ready ),
       .io_smi_req_valid( scr_conv_io_smi_req_valid ),
       .io_smi_req_bits_rw( scr_conv_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( scr_conv_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( scr_conv_io_smi_req_bits_data ),
       .io_smi_resp_ready( scr_conv_io_smi_resp_ready ),
       .io_smi_resp_valid( io_scr_resp_valid ),
       .io_smi_resp_bits( io_scr_resp_bits )
  );
endmodule

module SCRFile(input clk, input reset,
    output io_smi_req_ready,
    input  io_smi_req_valid,
    input  io_smi_req_bits_rw,
    input [5:0] io_smi_req_bits_addr,
    input [63:0] io_smi_req_bits_data,
    input  io_smi_resp_ready,
    output io_smi_resp_valid,
    output[63:0] io_smi_resp_bits,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    input [63:0] io_scr_rdata_1,
    input [63:0] io_scr_rdata_0,
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[63:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T8;
  wire[5:0] T9;
  reg [5:0] read_addr;
  wire[5:0] T135;
  wire[5:0] T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T13;
  wire T14;
  wire[63:0] T15;
  wire[63:0] T16;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T17;
  wire[63:0] T18;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T19;
  wire T20;
  wire T21;
  wire[63:0] T22;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T25;
  wire[63:0] T26;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T27;
  wire T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T31;
  wire[63:0] T32;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T41;
  wire[63:0] T42;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T43;
  wire T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T47;
  wire[63:0] T48;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T49;
  wire T50;
  wire T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T55;
  wire[63:0] T56;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T57;
  wire T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T61;
  wire[63:0] T62;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire[63:0] T72;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T73;
  wire[63:0] T74;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T75;
  wire T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T79;
  wire[63:0] T80;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T81;
  wire T82;
  wire T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T87;
  wire[63:0] T88;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T89;
  wire T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T93;
  wire[63:0] T94;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[63:0] T99;
  wire[63:0] T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T103;
  wire[63:0] T104;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T105;
  wire T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T109;
  wire[63:0] T110;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T111;
  wire T112;
  wire T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T117;
  wire[63:0] T118;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T119;
  wire T120;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T123;
  wire[63:0] T124;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  reg  resp_valid;
  wire T136;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    read_addr = {1{$random}};
    resp_valid = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_scr_wdata = io_smi_req_bits_data;
  assign io_scr_waddr = io_smi_req_bits_addr;
  assign io_scr_wen = T0;
  assign T0 = T1 & io_smi_req_bits_rw;
  assign T1 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_resp_bits = T2;
  assign T2 = T130 ? T68 : T3;
  assign T3 = T67 ? T37 : T4;
  assign T4 = T36 ? T22 : T5;
  assign T5 = T21 ? T15 : T6;
  assign T6 = T14 ? T12 : T7;
  assign T7 = T8 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = io_scr_rdata_0;
  assign scr_rdata_1 = io_scr_rdata_1;
  assign T8 = T9[1'h0];
  assign T9 = read_addr;
  assign T135 = reset ? 6'h0 : T10;
  assign T10 = T11 ? io_smi_req_bits_addr : read_addr;
  assign T11 = io_smi_req_ready & io_smi_req_valid;
  assign T12 = T13 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T13 = T9[1'h0];
  assign T14 = T9[1'h1];
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T17 = T9[1'h0];
  assign T18 = T19 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T19 = T9[1'h0];
  assign T20 = T9[1'h1];
  assign T21 = T9[2'h2];
  assign T22 = T35 ? T29 : T23;
  assign T23 = T28 ? T26 : T24;
  assign T24 = T25 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T25 = T9[1'h0];
  assign T26 = T27 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T27 = T9[1'h0];
  assign T28 = T9[1'h1];
  assign T29 = T34 ? T32 : T30;
  assign T30 = T31 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T31 = T9[1'h0];
  assign T32 = T33 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T33 = T9[1'h0];
  assign T34 = T9[1'h1];
  assign T35 = T9[2'h2];
  assign T36 = T9[2'h3];
  assign T37 = T66 ? T52 : T38;
  assign T38 = T51 ? T45 : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T41 = T9[1'h0];
  assign T42 = T43 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T43 = T9[1'h0];
  assign T44 = T9[1'h1];
  assign T45 = T50 ? T48 : T46;
  assign T46 = T47 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T47 = T9[1'h0];
  assign T48 = T49 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T49 = T9[1'h0];
  assign T50 = T9[1'h1];
  assign T51 = T9[2'h2];
  assign T52 = T65 ? T59 : T53;
  assign T53 = T58 ? T56 : T54;
  assign T54 = T55 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T55 = T9[1'h0];
  assign T56 = T57 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T57 = T9[1'h0];
  assign T58 = T9[1'h1];
  assign T59 = T64 ? T62 : T60;
  assign T60 = T61 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T61 = T9[1'h0];
  assign T62 = T63 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T63 = T9[1'h0];
  assign T64 = T9[1'h1];
  assign T65 = T9[2'h2];
  assign T66 = T9[2'h3];
  assign T67 = T9[3'h4];
  assign T68 = T129 ? T99 : T69;
  assign T69 = T98 ? T84 : T70;
  assign T70 = T83 ? T77 : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T73 = T9[1'h0];
  assign T74 = T75 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T75 = T9[1'h0];
  assign T76 = T9[1'h1];
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T79 = T9[1'h0];
  assign T80 = T81 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T81 = T9[1'h0];
  assign T82 = T9[1'h1];
  assign T83 = T9[2'h2];
  assign T84 = T97 ? T91 : T85;
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T87 = T9[1'h0];
  assign T88 = T89 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T89 = T9[1'h0];
  assign T90 = T9[1'h1];
  assign T91 = T96 ? T94 : T92;
  assign T92 = T93 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T93 = T9[1'h0];
  assign T94 = T95 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T95 = T9[1'h0];
  assign T96 = T9[1'h1];
  assign T97 = T9[2'h2];
  assign T98 = T9[2'h3];
  assign T99 = T128 ? T114 : T100;
  assign T100 = T113 ? T107 : T101;
  assign T101 = T106 ? T104 : T102;
  assign T102 = T103 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T103 = T9[1'h0];
  assign T104 = T105 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T105 = T9[1'h0];
  assign T106 = T9[1'h1];
  assign T107 = T112 ? T110 : T108;
  assign T108 = T109 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T109 = T9[1'h0];
  assign T110 = T111 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T111 = T9[1'h0];
  assign T112 = T9[1'h1];
  assign T113 = T9[2'h2];
  assign T114 = T127 ? T121 : T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T117 = T9[1'h0];
  assign T118 = T119 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T119 = T9[1'h0];
  assign T120 = T9[1'h1];
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T123 = T9[1'h0];
  assign T124 = T125 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T125 = T9[1'h0];
  assign T126 = T9[1'h1];
  assign T127 = T9[2'h2];
  assign T128 = T9[2'h3];
  assign T129 = T9[3'h4];
  assign T130 = T9[3'h5];
  assign io_smi_resp_valid = resp_valid;
  assign T136 = reset ? 1'h0 : T131;
  assign T131 = T133 ? 1'h0 : T132;
  assign T132 = T11 ? 1'h1 : resp_valid;
  assign T133 = io_smi_resp_ready & io_smi_resp_valid;
  assign io_smi_req_ready = T134;
  assign T134 = resp_valid ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      read_addr <= 6'h0;
    end else if(T11) begin
      read_addr <= io_smi_req_bits_addr;
    end
    if(reset) begin
      resp_valid <= 1'h0;
    end else if(T133) begin
      resp_valid <= 1'h0;
    end else if(T11) begin
      resp_valid <= 1'h1;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_len,
    input [2:0] io_enq_bits_size,
    input [1:0] io_enq_bits_burst,
    input  io_enq_bits_lock,
    input [3:0] io_enq_bits_cache,
    input [2:0] io_enq_bits_prot,
    input [3:0] io_enq_bits_qos,
    input [3:0] io_enq_bits_region,
    input [5:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_len,
    output[2:0] io_deq_bits_size,
    output[1:0] io_deq_bits_burst,
    output io_deq_bits_lock,
    output[3:0] io_deq_bits_cache,
    output[2:0] io_deq_bits_prot,
    output[3:0] io_deq_bits_qos,
    output[3:0] io_deq_bits_region,
    output[5:0] io_deq_bits_id,
    output io_deq_bits_user,
    output io_count
);

  wire T29;
  wire[1:0] T0;
  reg  full;
  wire T30;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire T3;
  wire[67:0] T4;
  reg [67:0] ram [0:0];
  wire[67:0] T5;
  wire[67:0] T6;
  wire[67:0] T7;
  wire[21:0] T8;
  wire[10:0] T9;
  wire[6:0] T10;
  wire[10:0] T11;
  wire[6:0] T12;
  wire[45:0] T13;
  wire[5:0] T14;
  wire[2:0] T15;
  wire[39:0] T16;
  wire[5:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[2:0] T24;
  wire[7:0] T25;
  wire[31:0] T26;
  wire T27;
  wire empty;
  wire T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T29;
  assign T29 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T30 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_user = T3;
  assign T3 = T4[1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T13, T8};
  assign T8 = {T11, T9};
  assign T9 = {io_enq_bits_region, T10};
  assign T10 = {io_enq_bits_id, io_enq_bits_user};
  assign T11 = {io_enq_bits_cache, T12};
  assign T12 = {io_enq_bits_prot, io_enq_bits_qos};
  assign T13 = {T16, T14};
  assign T14 = {io_enq_bits_size, T15};
  assign T15 = {io_enq_bits_burst, io_enq_bits_lock};
  assign T16 = {io_enq_bits_addr, io_enq_bits_len};
  assign io_deq_bits_id = T17;
  assign T17 = T4[3'h6:1'h1];
  assign io_deq_bits_region = T18;
  assign T18 = T4[4'ha:3'h7];
  assign io_deq_bits_qos = T19;
  assign T19 = T4[4'he:4'hb];
  assign io_deq_bits_prot = T20;
  assign T20 = T4[5'h11:4'hf];
  assign io_deq_bits_cache = T21;
  assign T21 = T4[5'h15:5'h12];
  assign io_deq_bits_lock = T22;
  assign T22 = T4[5'h16];
  assign io_deq_bits_burst = T23;
  assign T23 = T4[5'h18:5'h17];
  assign io_deq_bits_size = T24;
  assign T24 = T4[5'h1b:5'h19];
  assign io_deq_bits_len = T25;
  assign T25 = T4[6'h23:5'h1c];
  assign io_deq_bits_addr = T26;
  assign T26 = T4[7'h43:6'h24];
  assign io_deq_valid = T27;
  assign T27 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module NastiROM(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [5:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    //output[1:0] io_b_bits_resp
    //output[5:0] io_b_bits_id
    //output io_b_bits_user
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [5:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[5:0] io_r_bits_id,
    output io_r_bits_user
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  reg  T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[5:0] T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] rdata;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[63:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire[63:0] T18;
  wire[31:0] T19;
  wire[31:0] T20;
  reg [63:0] rdata_word;
  wire[6:0] T22;
  wire[31:0] T23;
  wire T24;
  wire[31:0] T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[31:0] T52;
  wire T28;
  wire T29;
  wire T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire T33;
  wire[1:0] T34;
  wire[15:0] T35;
  wire T36;
  wire[47:0] T37;
  wire[47:0] T38;
  wire[47:0] T39;
  wire[47:0] T53;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire[55:0] T45;
  wire[55:0] T46;
  wire[55:0] T47;
  wire[55:0] T54;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[31:0] Queue_io_deq_bits_addr;
  wire[7:0] Queue_io_deq_bits_len;
  wire[2:0] Queue_io_deq_bits_size;
  wire[5:0] Queue_io_deq_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T4 = 1'b0;
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_b_bits_user = {1{$random}};
//  assign io_b_bits_id = {1{$random}};
//  assign io_b_bits_resp = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_aw_valid | io_w_valid;
  assign T5 = T6 | reset;
  assign T6 = T8 | T7;
  assign T7 = Queue_io_deq_bits_len == 8'h0;
  assign T8 = Queue_io_deq_valid ^ 1'h1;
  assign io_r_bits_user = T9;
  assign T9 = 1'h0;
  assign io_r_bits_id = T10;
  assign T10 = Queue_io_deq_bits_id;
  assign io_r_bits_last = T11;
  assign T11 = 1'h1;
  assign io_r_bits_data = T12;
  assign T12 = rdata;
  assign rdata = {T45, T13};
  assign T13 = T44 ? T43 : T14;
  assign T14 = T15[3'h7:1'h0];
  assign T15 = {T37, T16};
  assign T16 = T36 ? T35 : T17;
  assign T17 = T18[4'hf:1'h0];
  assign T18 = {T25, T19};
  assign T19 = T24 ? T23 : T20;
  assign T20 = rdata_word[5'h1f:1'h0];
  always @(*) case (T22)
    0: rdata_word = 64'hb020000edfe0dd0;
    1: rdata_word = 64'hc001000038000000;
    2: rdata_word = 64'h1100000028000000;
    3: rdata_word = 64'h10000000;
    4: rdata_word = 64'h880100004b000000;
    5: rdata_word = 64'h0;
    6: rdata_word = 64'h0;
    7: rdata_word = 64'h1000000;
    8: rdata_word = 64'h400000003000000;
    9: rdata_word = 64'h200000000000000;
    10: rdata_word = 64'h400000003000000;
    11: rdata_word = 64'h20000000f000000;
    12: rdata_word = 64'hc00000003000000;
    13: rdata_word = 64'h6b636f521b000000;
    14: rdata_word = 64'h706968432d7465;
    15: rdata_word = 64'h6f6d656d01000000;
    16: rdata_word = 64'h30407972;
    17: rdata_word = 64'h700000003000000;
    18: rdata_word = 64'h6f6d656d21000000;
    19: rdata_word = 64'h300000000007972;
    20: rdata_word = 64'h2d00000010000000;
    21: rdata_word = 64'h0;
    22: rdata_word = 64'h4000000000;
    23: rdata_word = 64'h100000002000000;
    24: rdata_word = 64'h73757063;
    25: rdata_word = 64'h400000003000000;
    26: rdata_word = 64'h200000000000000;
    27: rdata_word = 64'h400000003000000;
    28: rdata_word = 64'h20000000f000000;
    29: rdata_word = 64'h4075706301000000;
    30: rdata_word = 64'h3030303830303034;
    31: rdata_word = 64'h300000000000000;
    32: rdata_word = 64'h2100000004000000;
    33: rdata_word = 64'h300000000757063;
    34: rdata_word = 64'h3100000006000000;
    35: rdata_word = 64'h7663736972;
    36: rdata_word = 64'h500000003000000;
    37: rdata_word = 64'h343676723c000000;
    38: rdata_word = 64'h300000000000000;
    39: rdata_word = 64'h2d00000008000000;
    40: rdata_word = 64'h80004000000000;
    41: rdata_word = 64'h200000002000000;
    42: rdata_word = 64'h4072637301000000;
    43: rdata_word = 64'h3030303031303034;
    44: rdata_word = 64'h300000000000000;
    45: rdata_word = 64'h2100000004000000;
    46: rdata_word = 64'h300000000726373;
    47: rdata_word = 64'h3100000006000000;
    48: rdata_word = 64'h7663736972;
    49: rdata_word = 64'h400000003000000;
    50: rdata_word = 64'h300000040000000;
    51: rdata_word = 64'h1000000003000000;
    52: rdata_word = 64'h2d000000;
    53: rdata_word = 64'h140;
    54: rdata_word = 64'h200000000020000;
    55: rdata_word = 64'h900000002000000;
    56: rdata_word = 64'h7373657264646123;
    57: rdata_word = 64'h2300736c6c65632d;
    58: rdata_word = 64'h6c65632d657a6973;
    59: rdata_word = 64'h6c65646f6d00736c;
    60: rdata_word = 64'h5f65636976656400;
    61: rdata_word = 64'h6765720065707974;
    62: rdata_word = 64'h697461706d6f6300;
    63: rdata_word = 64'h61736900656c62;
    64: rdata_word = 64'h69746365746f7270;
    65: rdata_word = 64'h6e6f;
    66: rdata_word = 64'h0;
    default: begin
      rdata_word = 64'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      rdata_word = {2{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T22 = Queue_io_deq_bits_addr[4'h9:2'h3];
  assign T23 = rdata_word[6'h3f:6'h20];
  assign T24 = Queue_io_deq_bits_addr[2'h2];
  assign T25 = T33 ? T27 : T26;
  assign T26 = rdata_word[6'h3f:6'h20];
  assign T27 = 32'h0 - T52;
  assign T52 = {31'h0, T28};
  assign T28 = T30 & T29;
  assign T29 = T19[5'h1f];
  assign T30 = $signed(1'h0) <= $signed(T31);
  assign T31 = T32;
  assign T32 = {1'h1, Queue_io_deq_bits_size};
  assign T33 = T34 == 2'h2;
  assign T34 = T32[1'h1:1'h0];
  assign T35 = T18[5'h1f:5'h10];
  assign T36 = Queue_io_deq_bits_addr[1'h1];
  assign T37 = T42 ? T39 : T38;
  assign T38 = T18[6'h3f:5'h10];
  assign T39 = 48'h0 - T53;
  assign T53 = {47'h0, T40};
  assign T40 = T30 & T41;
  assign T41 = T16[4'hf];
  assign T42 = T34 == 2'h1;
  assign T43 = T15[4'hf:4'h8];
  assign T44 = Queue_io_deq_bits_addr[1'h0];
  assign T45 = T50 ? T47 : T46;
  assign T46 = T15[6'h3f:4'h8];
  assign T47 = 56'h0 - T54;
  assign T54 = {55'h0, T48};
  assign T48 = T30 & T49;
  assign T49 = T13[3'h7];
  assign T50 = T34 == 2'h0;
  assign io_r_bits_resp = T51;
  assign T51 = 2'h0;
  assign io_r_valid = Queue_io_deq_valid;
  assign io_ar_ready = Queue_io_enq_ready;
  assign io_b_valid = 1'h0;
  assign io_w_ready = 1'h0;
  assign io_aw_ready = 1'h0;
  Queue_7 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_ar_valid ),
       .io_enq_bits_addr( io_ar_bits_addr ),
       .io_enq_bits_len( io_ar_bits_len ),
       .io_enq_bits_size( io_ar_bits_size ),
       .io_enq_bits_burst( io_ar_bits_burst ),
       .io_enq_bits_lock( io_ar_bits_lock ),
       .io_enq_bits_cache( io_ar_bits_cache ),
       .io_enq_bits_prot( io_ar_bits_prot ),
       .io_enq_bits_qos( io_ar_bits_qos ),
       .io_enq_bits_region( io_ar_bits_region ),
       .io_enq_bits_id( io_ar_bits_id ),
       .io_enq_bits_user( io_ar_bits_user ),
       .io_deq_ready( io_r_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_io_deq_bits_len ),
       .io_deq_bits_size( Queue_io_deq_bits_size ),
       //.io_deq_bits_burst(  )
       //.io_deq_bits_lock(  )
       //.io_deq_bits_cache(  )
       //.io_deq_bits_prot(  )
       //.io_deq_bits_qos(  )
       //.io_deq_bits_region(  )
       .io_deq_bits_id( Queue_io_deq_bits_id )
       //.io_deq_bits_user(  )
       //.io_count(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T4 <= 1'b1;
  if(!T5 && T4 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't burst-read from NastiROM");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't write to NastiROM");
    $finish;
  end
// synthesis translate_on
`endif
  end
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [16:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[16:0] io_deq_bits,
    output io_count
);

  wire T7;
  wire[1:0] T0;
  reg  full;
  wire T8;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[16:0] T3;
  reg [16:0] ram [0:0];
  wire[16:0] T4;
  wire T5;
  wire empty;
  wire T6;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T7;
  assign T7 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T8 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits = T3;
  assign T3 = ram[1'h0];
  assign io_deq_valid = T5;
  assign T5 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T6;
  assign T6 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= io_enq_bits;
  end
endmodule

module SlowIO(input clk, input reset,
    output io_out_fast_ready,
    input  io_out_fast_valid,
    input [16:0] io_out_fast_bits,
    input  io_out_slow_ready,
    output io_out_slow_valid,
    output[16:0] io_out_slow_bits,
    input  io_in_fast_ready,
    output io_in_fast_valid,
    output[16:0] io_in_fast_bits,
    output io_in_slow_ready,
    input  io_in_slow_valid,
    input [16:0] io_in_slow_bits,
    output io_clk_slow,
    input  io_set_divisor_valid,
    input [31:0] io_set_divisor_bits,
    output[31:0] io_divisor
);

  wire T0;
  reg  out_slow_val;
  wire T26;
  wire T1;
  wire held;
  wire[8:0] T2;
  reg [8:0] hold;
  wire[8:0] T27;
  wire[8:0] T3;
  reg [8:0] h_shadow;
  wire[8:0] T28;
  wire[8:0] T4;
  wire[8:0] T5;
  wire[8:0] T6;
  wire falling;
  reg [8:0] divisor;
  wire[8:0] T29;
  wire[8:0] T7;
  reg [8:0] d_shadow;
  wire[8:0] T30;
  wire[8:0] T8;
  wire[8:0] T9;
  wire[8:0] T10;
  wire[8:0] T31;
  wire[7:0] T11;
  reg [8:0] count;
  wire[8:0] T12;
  wire[8:0] T13;
  wire T14;
  wire rising;
  wire[8:0] T32;
  wire[7:0] T15;
  wire T16;
  wire T17;
  wire T18;
  reg  in_slow_rdy;
  wire T33;
  wire T19;
  wire[31:0] T34;
  wire[24:0] T20;
  wire[24:0] T35;
  wire[24:0] T21;
  reg  myclock;
  wire T22;
  wire T23;
  reg [16:0] out_slow_bits;
  wire[16:0] T24;
  wire[16:0] T25;
  wire fromhost_q_io_enq_ready;
  wire fromhost_q_io_deq_valid;
  wire[16:0] fromhost_q_io_deq_bits;
  wire tohost_q_io_enq_ready;
  wire tohost_q_io_deq_valid;
  wire[16:0] tohost_q_io_deq_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_slow_val = {1{$random}};
    hold = {1{$random}};
    h_shadow = {1{$random}};
    divisor = {1{$random}};
    d_shadow = {1{$random}};
    count = {1{$random}};
    in_slow_rdy = {1{$random}};
    myclock = {1{$random}};
    out_slow_bits = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T14 & out_slow_val;
  assign T26 = reset ? 1'h0 : T1;
  assign T1 = held ? tohost_q_io_deq_valid : out_slow_val;
  assign held = count == T2;
  assign T2 = T31 + hold;
  assign T27 = reset ? 9'h7f : T3;
  assign T3 = falling ? h_shadow : hold;
  assign T28 = reset ? 9'h7f : T4;
  assign T4 = io_set_divisor_valid ? T5 : h_shadow;
  assign T5 = T6;
  assign T6 = io_set_divisor_bits[5'h18:5'h10];
  assign falling = count == divisor;
  assign T29 = reset ? 9'h1ff : T7;
  assign T7 = falling ? d_shadow : divisor;
  assign T30 = reset ? 9'h1ff : T8;
  assign T8 = io_set_divisor_valid ? T9 : d_shadow;
  assign T9 = T10;
  assign T10 = io_set_divisor_bits[4'h8:1'h0];
  assign T31 = {1'h0, T11};
  assign T11 = divisor >> 1'h1;
  assign T12 = falling ? 9'h0 : T13;
  assign T13 = count + 9'h1;
  assign T14 = rising & io_out_slow_ready;
  assign rising = count == T32;
  assign T32 = {1'h0, T15};
  assign T15 = divisor >> 1'h1;
  assign T16 = rising & T17;
  assign T17 = T18 | reset;
  assign T18 = io_in_slow_valid & in_slow_rdy;
  assign T33 = reset ? 1'h0 : T19;
  assign T19 = held ? fromhost_q_io_enq_ready : in_slow_rdy;
  assign io_divisor = T34;
  assign T34 = {7'h0, T20};
  assign T20 = T21 | T35;
  assign T35 = {16'h0, divisor};
  assign T21 = hold << 5'h10;
  assign io_clk_slow = myclock;
  assign T22 = rising ? 1'h1 : T23;
  assign T23 = falling ? 1'h0 : myclock;
  assign io_in_slow_ready = in_slow_rdy;
  assign io_in_fast_bits = fromhost_q_io_deq_bits;
  assign io_in_fast_valid = fromhost_q_io_deq_valid;
  assign io_out_slow_bits = out_slow_bits;
  assign T24 = held ? T25 : out_slow_bits;
  assign T25 = reset ? fromhost_q_io_deq_bits : tohost_q_io_deq_bits;
  assign io_out_slow_valid = out_slow_val;
  assign io_out_fast_ready = tohost_q_io_enq_ready;
  Queue_8 fromhost_q(.clk(clk), .reset(reset),
       .io_enq_ready( fromhost_q_io_enq_ready ),
       .io_enq_valid( T16 ),
       .io_enq_bits( io_in_slow_bits ),
       .io_deq_ready( io_in_fast_ready ),
       .io_deq_valid( fromhost_q_io_deq_valid ),
       .io_deq_bits( fromhost_q_io_deq_bits )
       //.io_count(  )
  );
  Queue_8 tohost_q(.clk(clk), .reset(reset),
       .io_enq_ready( tohost_q_io_enq_ready ),
       .io_enq_valid( io_out_fast_valid ),
       .io_enq_bits( io_out_fast_bits ),
       .io_deq_ready( T0 ),
       .io_deq_valid( tohost_q_io_deq_valid ),
       .io_deq_bits( tohost_q_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      out_slow_val <= 1'h0;
    end else if(held) begin
      out_slow_val <= tohost_q_io_deq_valid;
    end
    if(reset) begin
      hold <= 9'h7f;
    end else if(falling) begin
      hold <= h_shadow;
    end
    if(reset) begin
      h_shadow <= 9'h7f;
    end else if(io_set_divisor_valid) begin
      h_shadow <= T5;
    end
    if(reset) begin
      divisor <= 9'h1ff;
    end else if(falling) begin
      divisor <= d_shadow;
    end
    if(reset) begin
      d_shadow <= 9'h1ff;
    end else if(io_set_divisor_valid) begin
      d_shadow <= T9;
    end
    if(falling) begin
      count <= 9'h0;
    end else begin
      count <= T13;
    end
    if(reset) begin
      in_slow_rdy <= 1'h0;
    end else if(held) begin
      in_slow_rdy <= fromhost_q_io_enq_ready;
    end
    if(rising) begin
      myclock <= 1'h1;
    end else if(falling) begin
      myclock <= 1'h0;
    end
    if(held) begin
      out_slow_bits <= T25;
    end
  end
endmodule

module Uncore(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[5:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [5:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[5:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [5:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [5:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[5:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [5:0] io_tiles_cached_0_release_bits_client_xact_id,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [5:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[5:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[3:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_0_reset,
    output io_htif_0_id,
    input  io_htif_0_csr_req_ready,
    output io_htif_0_csr_req_valid,
    output io_htif_0_csr_req_bits_rw,
    output[11:0] io_htif_0_csr_req_bits_addr,
    output[63:0] io_htif_0_csr_req_bits_data,
    output io_htif_0_csr_resp_ready,
    input  io_htif_0_csr_resp_valid,
    input [63:0] io_htif_0_csr_resp_bits,
    input  io_htif_0_debug_stats_csr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    output io_mem_backup_ctrl_out_valid
    //input  io_mmio_aw_ready
    //output io_mmio_aw_valid
    //output[31:0] io_mmio_aw_bits_addr
    //output[7:0] io_mmio_aw_bits_len
    //output[2:0] io_mmio_aw_bits_size
    //output[1:0] io_mmio_aw_bits_burst
    //output io_mmio_aw_bits_lock
    //output[3:0] io_mmio_aw_bits_cache
    //output[2:0] io_mmio_aw_bits_prot
    //output[3:0] io_mmio_aw_bits_qos
    //output[3:0] io_mmio_aw_bits_region
    //output[5:0] io_mmio_aw_bits_id
    //output io_mmio_aw_bits_user
    //input  io_mmio_w_ready
    //output io_mmio_w_valid
    //output[63:0] io_mmio_w_bits_data
    //output io_mmio_w_bits_last
    //output[7:0] io_mmio_w_bits_strb
    //output io_mmio_w_bits_user
    //output io_mmio_b_ready
    //input  io_mmio_b_valid
    //input [1:0] io_mmio_b_bits_resp
    //input [5:0] io_mmio_b_bits_id
    //input  io_mmio_b_bits_user
    //input  io_mmio_ar_ready
    //output io_mmio_ar_valid
    //output[31:0] io_mmio_ar_bits_addr
    //output[7:0] io_mmio_ar_bits_len
    //output[2:0] io_mmio_ar_bits_size
    //output[1:0] io_mmio_ar_bits_burst
    //output io_mmio_ar_bits_lock
    //output[3:0] io_mmio_ar_bits_cache
    //output[2:0] io_mmio_ar_bits_prot
    //output[3:0] io_mmio_ar_bits_qos
    //output[3:0] io_mmio_ar_bits_region
    //output[5:0] io_mmio_ar_bits_id
    //output io_mmio_ar_bits_user
    //output io_mmio_r_ready
    //input  io_mmio_r_valid
    //input [1:0] io_mmio_r_bits_resp
    //input [63:0] io_mmio_r_bits_data
    //input  io_mmio_r_bits_last
    //input [5:0] io_mmio_r_bits_id
    //input  io_mmio_r_bits_user
);

  wire[31:0] T33;
  wire T0;
  wire T1;
  wire[16:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[16:0] T9;
  wire[15:0] T10;
  wire T11;
  wire[63:0] T12;
  reg  memory_channel_mux_select;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[63:0] T34;
  wire[15:0] T35;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[15:0] T36;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[15:0] T37;
  wire T27;
  wire T28;
  reg  R29;
  wire T30;
  wire T31;
  reg  R32;
  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_csr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_id;
  wire htif_io_cpu_0_csr_req_valid;
  wire htif_io_cpu_0_csr_req_bits_rw;
  wire[11:0] htif_io_cpu_0_csr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_csr_req_bits_data;
  wire htif_io_cpu_0_csr_resp_ready;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_addr_block;
  wire[5:0] htif_io_mem_acquire_bits_client_xact_id;
  wire[1:0] htif_io_mem_acquire_bits_addr_beat;
  wire htif_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] htif_io_mem_acquire_bits_a_type;
  wire[16:0] htif_io_mem_acquire_bits_union;
  wire[127:0] htif_io_mem_acquire_bits_data;
  wire htif_io_mem_grant_ready;
  wire htif_io_scr_req_valid;
  wire htif_io_scr_req_bits_rw;
  wire[5:0] htif_io_scr_req_bits_addr;
  wire[63:0] htif_io_scr_req_bits_data;
  wire htif_io_scr_resp_ready;
  wire scrFile_io_smi_req_ready;
  wire scrFile_io_smi_resp_valid;
  wire[63:0] scrFile_io_smi_resp_bits;
  wire scrFile_io_scr_wen;
  wire[5:0] scrFile_io_scr_waddr;
  wire[63:0] scrFile_io_scr_wdata;
  wire SmiArbiter_io_in_1_req_ready;
  wire SmiArbiter_io_in_1_resp_valid;
  wire[63:0] SmiArbiter_io_in_1_resp_bits;
  wire SmiArbiter_io_in_0_req_ready;
  wire SmiArbiter_io_in_0_resp_valid;
  wire[63:0] SmiArbiter_io_in_0_resp_bits;
  wire SmiArbiter_io_out_req_valid;
  wire SmiArbiter_io_out_req_bits_rw;
  wire[11:0] SmiArbiter_io_out_req_bits_addr;
  wire[63:0] SmiArbiter_io_out_req_bits_data;
  wire SmiArbiter_io_out_resp_ready;
  wire scrArb_io_in_1_req_ready;
  wire scrArb_io_in_1_resp_valid;
  wire[63:0] scrArb_io_in_1_resp_bits;
  wire scrArb_io_in_0_req_ready;
  wire scrArb_io_in_0_resp_valid;
  wire[63:0] scrArb_io_in_0_resp_bits;
  wire scrArb_io_out_req_valid;
  wire scrArb_io_out_req_bits_rw;
  wire[5:0] scrArb_io_out_req_bits_addr;
  wire[63:0] scrArb_io_out_req_bits_data;
  wire scrArb_io_out_resp_ready;
  wire deviceTree_io_aw_ready;
  wire deviceTree_io_w_ready;
  wire deviceTree_io_b_valid;
  wire deviceTree_io_ar_ready;
  wire deviceTree_io_r_valid;
  wire[1:0] deviceTree_io_r_bits_resp;
  wire[63:0] deviceTree_io_r_bits_data;
  wire deviceTree_io_r_bits_last;
  wire[5:0] deviceTree_io_r_bits_id;
  wire deviceTree_io_r_bits_user;
  wire SlowIO_io_out_fast_ready;
  wire SlowIO_io_out_slow_valid;
  wire[16:0] SlowIO_io_out_slow_bits;
  wire SlowIO_io_in_fast_valid;
  wire[16:0] SlowIO_io_in_fast_bits;
  wire SlowIO_io_in_slow_ready;
  wire SlowIO_io_clk_slow;
  wire[31:0] SlowIO_io_divisor;
  wire outmemsys_io_tiles_cached_0_acquire_ready;
  wire outmemsys_io_tiles_cached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire[5:0] outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire outmemsys_io_tiles_cached_0_probe_valid;
  wire[25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire outmemsys_io_tiles_cached_0_release_ready;
  wire outmemsys_io_tiles_uncached_0_acquire_ready;
  wire outmemsys_io_tiles_uncached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[5:0] outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire outmemsys_io_htif_uncached_acquire_ready;
  wire outmemsys_io_htif_uncached_grant_valid;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_addr_beat;
  wire[5:0] outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  wire outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_g_type;
  wire[127:0] outmemsys_io_htif_uncached_grant_bits_data;
  wire outmemsys_io_mem_0_aw_valid;
  wire[31:0] outmemsys_io_mem_0_aw_bits_addr;
  wire[7:0] outmemsys_io_mem_0_aw_bits_len;
  wire[2:0] outmemsys_io_mem_0_aw_bits_size;
  wire[1:0] outmemsys_io_mem_0_aw_bits_burst;
  wire outmemsys_io_mem_0_aw_bits_lock;
  wire[3:0] outmemsys_io_mem_0_aw_bits_cache;
  wire[2:0] outmemsys_io_mem_0_aw_bits_prot;
  wire[3:0] outmemsys_io_mem_0_aw_bits_qos;
  wire[3:0] outmemsys_io_mem_0_aw_bits_region;
  wire[5:0] outmemsys_io_mem_0_aw_bits_id;
  wire outmemsys_io_mem_0_aw_bits_user;
  wire outmemsys_io_mem_0_w_valid;
  wire[63:0] outmemsys_io_mem_0_w_bits_data;
  wire outmemsys_io_mem_0_w_bits_last;
  wire[7:0] outmemsys_io_mem_0_w_bits_strb;
  wire outmemsys_io_mem_0_w_bits_user;
  wire outmemsys_io_mem_0_b_ready;
  wire outmemsys_io_mem_0_ar_valid;
  wire[31:0] outmemsys_io_mem_0_ar_bits_addr;
  wire[7:0] outmemsys_io_mem_0_ar_bits_len;
  wire[2:0] outmemsys_io_mem_0_ar_bits_size;
  wire[1:0] outmemsys_io_mem_0_ar_bits_burst;
  wire outmemsys_io_mem_0_ar_bits_lock;
  wire[3:0] outmemsys_io_mem_0_ar_bits_cache;
  wire[2:0] outmemsys_io_mem_0_ar_bits_prot;
  wire[3:0] outmemsys_io_mem_0_ar_bits_qos;
  wire[3:0] outmemsys_io_mem_0_ar_bits_region;
  wire[5:0] outmemsys_io_mem_0_ar_bits_id;
  wire outmemsys_io_mem_0_ar_bits_user;
  wire outmemsys_io_mem_0_r_ready;
  wire outmemsys_io_mem_backup_req_valid;
  wire[15:0] outmemsys_io_mem_backup_req_bits;
  wire outmemsys_io_csr_0_req_valid;
  wire outmemsys_io_csr_0_req_bits_rw;
  wire[11:0] outmemsys_io_csr_0_req_bits_addr;
  wire[63:0] outmemsys_io_csr_0_req_bits_data;
  wire outmemsys_io_csr_0_resp_ready;
  wire outmemsys_io_scr_req_valid;
  wire outmemsys_io_scr_req_bits_rw;
  wire[5:0] outmemsys_io_scr_req_bits_addr;
  wire[63:0] outmemsys_io_scr_req_bits_data;
  wire outmemsys_io_scr_resp_ready;
  wire outmemsys_io_deviceTree_aw_valid;
  wire[31:0] outmemsys_io_deviceTree_aw_bits_addr;
  wire[7:0] outmemsys_io_deviceTree_aw_bits_len;
  wire[2:0] outmemsys_io_deviceTree_aw_bits_size;
  wire[1:0] outmemsys_io_deviceTree_aw_bits_burst;
  wire outmemsys_io_deviceTree_aw_bits_lock;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_cache;
  wire[2:0] outmemsys_io_deviceTree_aw_bits_prot;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_qos;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_region;
  wire[5:0] outmemsys_io_deviceTree_aw_bits_id;
  wire outmemsys_io_deviceTree_aw_bits_user;
  wire outmemsys_io_deviceTree_w_valid;
  wire[63:0] outmemsys_io_deviceTree_w_bits_data;
  wire outmemsys_io_deviceTree_w_bits_last;
  wire[7:0] outmemsys_io_deviceTree_w_bits_strb;
  wire outmemsys_io_deviceTree_w_bits_user;
  wire outmemsys_io_deviceTree_b_ready;
  wire outmemsys_io_deviceTree_ar_valid;
  wire[31:0] outmemsys_io_deviceTree_ar_bits_addr;
  wire[7:0] outmemsys_io_deviceTree_ar_bits_len;
  wire[2:0] outmemsys_io_deviceTree_ar_bits_size;
  wire[1:0] outmemsys_io_deviceTree_ar_bits_burst;
  wire outmemsys_io_deviceTree_ar_bits_lock;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_cache;
  wire[2:0] outmemsys_io_deviceTree_ar_bits_prot;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_qos;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_region;
  wire[5:0] outmemsys_io_deviceTree_ar_bits_id;
  wire outmemsys_io_deviceTree_ar_bits_user;
  wire outmemsys_io_deviceTree_r_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    memory_channel_mux_select = {1{$random}};
    R29 = {1{$random}};
    R32 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mmio_r_ready = {1{$random}};
//  assign io_mmio_ar_bits_user = {1{$random}};
//  assign io_mmio_ar_bits_id = {1{$random}};
//  assign io_mmio_ar_bits_region = {1{$random}};
//  assign io_mmio_ar_bits_qos = {1{$random}};
//  assign io_mmio_ar_bits_prot = {1{$random}};
//  assign io_mmio_ar_bits_cache = {1{$random}};
//  assign io_mmio_ar_bits_lock = {1{$random}};
//  assign io_mmio_ar_bits_burst = {1{$random}};
//  assign io_mmio_ar_bits_size = {1{$random}};
//  assign io_mmio_ar_bits_len = {1{$random}};
//  assign io_mmio_ar_bits_addr = {1{$random}};
//  assign io_mmio_ar_valid = {1{$random}};
//  assign io_mmio_b_ready = {1{$random}};
//  assign io_mmio_w_bits_user = {1{$random}};
//  assign io_mmio_w_bits_strb = {1{$random}};
//  assign io_mmio_w_bits_last = {1{$random}};
//  assign io_mmio_w_bits_data = {2{$random}};
//  assign io_mmio_w_valid = {1{$random}};
//  assign io_mmio_aw_bits_user = {1{$random}};
//  assign io_mmio_aw_bits_id = {1{$random}};
//  assign io_mmio_aw_bits_region = {1{$random}};
//  assign io_mmio_aw_bits_qos = {1{$random}};
//  assign io_mmio_aw_bits_prot = {1{$random}};
//  assign io_mmio_aw_bits_cache = {1{$random}};
//  assign io_mmio_aw_bits_lock = {1{$random}};
//  assign io_mmio_aw_bits_burst = {1{$random}};
//  assign io_mmio_aw_bits_size = {1{$random}};
//  assign io_mmio_aw_bits_len = {1{$random}};
//  assign io_mmio_aw_bits_addr = {1{$random}};
//  assign io_mmio_aw_valid = {1{$random}};
// synthesis translate_on
`endif
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign T33 = scrFile_io_scr_wdata[5'h1f:1'h0];
  assign T0 = scrFile_io_scr_wen & T1;
  assign T1 = scrFile_io_scr_waddr == 6'h3f;
  assign T2 = {T3, io_host_in_bits};
  assign T3 = io_mem_backup_ctrl_en & io_mem_backup_ctrl_in_valid;
  assign T4 = T3 | io_host_in_valid;
  assign T5 = T6 ? 1'h1 : htif_io_host_in_ready;
  assign T6 = SlowIO_io_in_fast_bits[5'h10];
  assign T7 = T8 ? io_host_out_ready : io_mem_backup_ctrl_out_ready;
  assign T8 = SlowIO_io_out_slow_bits[5'h10];
  assign T9 = {htif_io_host_out_valid, T10};
  assign T10 = htif_io_host_out_valid ? htif_io_host_out_bits : outmemsys_io_mem_backup_req_bits;
  assign T11 = htif_io_host_out_valid | outmemsys_io_mem_backup_req_valid;
  assign T12 = {63'h0, memory_channel_mux_select};
  assign T13 = T15 ? T14 : memory_channel_mux_select;
  assign T14 = scrFile_io_scr_wdata[1'h0];
  assign T15 = scrFile_io_scr_wen & T16;
  assign T16 = scrFile_io_scr_waddr == 6'h2;
  assign T34 = {32'h0, SlowIO_io_divisor};
  assign T35 = SlowIO_io_in_fast_bits[4'hf:1'h0];
  assign T17 = SlowIO_io_in_fast_valid & T18;
  assign T18 = SlowIO_io_in_fast_bits[5'h10];
  assign T19 = SlowIO_io_out_fast_ready & T20;
  assign T20 = htif_io_host_out_valid ^ 1'h1;
  assign T36 = SlowIO_io_in_fast_bits[4'hf:1'h0];
  assign T21 = SlowIO_io_in_fast_valid & T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = SlowIO_io_in_fast_bits[5'h10];
  assign io_mem_backup_ctrl_out_valid = T24;
  assign T24 = SlowIO_io_out_slow_valid & T25;
  assign T25 = T26 ^ 1'h1;
  assign T26 = SlowIO_io_out_slow_bits[5'h10];
  assign io_htif_0_csr_resp_ready = SmiArbiter_io_out_resp_ready;
  assign io_htif_0_csr_req_bits_data = SmiArbiter_io_out_req_bits_data;
  assign io_htif_0_csr_req_bits_addr = SmiArbiter_io_out_req_bits_addr;
  assign io_htif_0_csr_req_bits_rw = SmiArbiter_io_out_req_bits_rw;
  assign io_htif_0_csr_req_valid = SmiArbiter_io_out_req_valid;
  assign io_htif_0_id = htif_io_cpu_0_id;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_mem_0_r_ready = outmemsys_io_mem_0_r_ready;
  assign io_mem_0_ar_bits_user = outmemsys_io_mem_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = outmemsys_io_mem_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = outmemsys_io_mem_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = outmemsys_io_mem_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = outmemsys_io_mem_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = outmemsys_io_mem_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = outmemsys_io_mem_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = outmemsys_io_mem_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = outmemsys_io_mem_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = outmemsys_io_mem_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = outmemsys_io_mem_0_ar_bits_addr;
  assign io_mem_0_ar_valid = outmemsys_io_mem_0_ar_valid;
  assign io_mem_0_b_ready = outmemsys_io_mem_0_b_ready;
  assign io_mem_0_w_bits_user = outmemsys_io_mem_0_w_bits_user;
  assign io_mem_0_w_bits_strb = outmemsys_io_mem_0_w_bits_strb;
  assign io_mem_0_w_bits_last = outmemsys_io_mem_0_w_bits_last;
  assign io_mem_0_w_bits_data = outmemsys_io_mem_0_w_bits_data;
  assign io_mem_0_w_valid = outmemsys_io_mem_0_w_valid;
  assign io_mem_0_aw_bits_user = outmemsys_io_mem_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = outmemsys_io_mem_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = outmemsys_io_mem_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = outmemsys_io_mem_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = outmemsys_io_mem_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = outmemsys_io_mem_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = outmemsys_io_mem_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = outmemsys_io_mem_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = outmemsys_io_mem_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = outmemsys_io_mem_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = outmemsys_io_mem_0_aw_bits_addr;
  assign io_mem_0_aw_valid = outmemsys_io_mem_0_aw_valid;
  assign io_host_debug_stats_csr = htif_io_host_debug_stats_csr;
  assign io_host_out_bits = T37;
  assign T37 = SlowIO_io_out_slow_bits[4'hf:1'h0];
  assign io_host_out_valid = T27;
  assign T27 = SlowIO_io_out_slow_valid & T28;
  assign T28 = SlowIO_io_out_slow_bits[5'h10];
  assign io_host_in_ready = SlowIO_io_in_slow_ready;
  assign io_host_clk_edge = R29;
  assign T30 = io_host_clk & T31;
  assign T31 = R32 ^ 1'h1;
  assign io_host_clk = SlowIO_io_clk_slow;
  Htif htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( T21 ),
       .io_host_in_bits( T36 ),
       .io_host_out_ready( SlowIO_io_out_fast_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_csr( htif_io_host_debug_stats_csr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       .io_cpu_0_id( htif_io_cpu_0_id ),
       .io_cpu_0_csr_req_ready( SmiArbiter_io_in_0_req_ready ),
       .io_cpu_0_csr_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_cpu_0_csr_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_cpu_0_csr_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_cpu_0_csr_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_cpu_0_csr_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_cpu_0_csr_resp_valid( SmiArbiter_io_in_0_resp_valid ),
       .io_cpu_0_csr_resp_bits( SmiArbiter_io_in_0_resp_bits ),
       .io_cpu_0_debug_stats_csr( io_htif_0_debug_stats_csr ),
       .io_mem_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_mem_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_mem_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_scr_req_ready( scrArb_io_in_0_req_ready ),
       .io_scr_req_valid( htif_io_scr_req_valid ),
       .io_scr_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( htif_io_scr_req_bits_data ),
       .io_scr_resp_ready( htif_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_0_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign htif.io_cpu_0_id = {1{$random}};
// synthesis translate_on
`endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_cached_0_acquire_ready( outmemsys_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( outmemsys_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( outmemsys_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( outmemsys_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( outmemsys_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( outmemsys_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( outmemsys_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( outmemsys_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( outmemsys_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( outmemsys_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( outmemsys_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( outmemsys_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( outmemsys_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( outmemsys_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( outmemsys_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_uncached_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_htif_uncached_acquire_valid( htif_io_mem_acquire_valid ),
       .io_htif_uncached_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_htif_uncached_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_htif_uncached_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_htif_uncached_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_htif_uncached_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_htif_uncached_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_htif_uncached_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_htif_uncached_grant_ready( htif_io_mem_grant_ready ),
       .io_htif_uncached_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_htif_uncached_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_htif_uncached_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_htif_uncached_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_htif_uncached_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_htif_uncached_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_htif_uncached_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_incoherent_0( htif_io_cpu_0_reset ),
       .io_mem_0_aw_ready( io_mem_0_aw_ready ),
       .io_mem_0_aw_valid( outmemsys_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( outmemsys_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( outmemsys_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( outmemsys_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( outmemsys_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( outmemsys_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( outmemsys_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( outmemsys_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( outmemsys_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( outmemsys_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( outmemsys_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( outmemsys_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( io_mem_0_w_ready ),
       .io_mem_0_w_valid( outmemsys_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( outmemsys_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( outmemsys_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( outmemsys_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( outmemsys_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( outmemsys_io_mem_0_b_ready ),
       .io_mem_0_b_valid( io_mem_0_b_valid ),
       .io_mem_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_mem_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_mem_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_mem_0_ar_ready( io_mem_0_ar_ready ),
       .io_mem_0_ar_valid( outmemsys_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( outmemsys_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( outmemsys_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( outmemsys_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( outmemsys_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( outmemsys_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( outmemsys_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( outmemsys_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( outmemsys_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( outmemsys_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( outmemsys_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( outmemsys_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( outmemsys_io_mem_0_r_ready ),
       .io_mem_0_r_valid( io_mem_0_r_valid ),
       .io_mem_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_mem_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_mem_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_mem_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_mem_0_r_bits_user( io_mem_0_r_bits_user ),
       .io_mem_backup_req_ready( T19 ),
       .io_mem_backup_req_valid( outmemsys_io_mem_backup_req_valid ),
       .io_mem_backup_req_bits( outmemsys_io_mem_backup_req_bits ),
       .io_mem_backup_resp_valid( T17 ),
       .io_mem_backup_resp_bits( T35 ),
       .io_mem_backup_en( io_mem_backup_ctrl_en ),
       .io_memory_channel_mux_select( memory_channel_mux_select ),
       .io_csr_0_req_ready( SmiArbiter_io_in_1_req_ready ),
       .io_csr_0_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_csr_0_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_csr_0_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_csr_0_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_csr_0_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_csr_0_resp_valid( SmiArbiter_io_in_1_resp_valid ),
       .io_csr_0_resp_bits( SmiArbiter_io_in_1_resp_bits ),
       .io_scr_req_ready( scrArb_io_in_1_req_ready ),
       .io_scr_req_valid( outmemsys_io_scr_req_valid ),
       .io_scr_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_scr_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_deviceTree_aw_ready( deviceTree_io_aw_ready ),
       .io_deviceTree_aw_valid( outmemsys_io_deviceTree_aw_valid ),
       .io_deviceTree_aw_bits_addr( outmemsys_io_deviceTree_aw_bits_addr ),
       .io_deviceTree_aw_bits_len( outmemsys_io_deviceTree_aw_bits_len ),
       .io_deviceTree_aw_bits_size( outmemsys_io_deviceTree_aw_bits_size ),
       .io_deviceTree_aw_bits_burst( outmemsys_io_deviceTree_aw_bits_burst ),
       .io_deviceTree_aw_bits_lock( outmemsys_io_deviceTree_aw_bits_lock ),
       .io_deviceTree_aw_bits_cache( outmemsys_io_deviceTree_aw_bits_cache ),
       .io_deviceTree_aw_bits_prot( outmemsys_io_deviceTree_aw_bits_prot ),
       .io_deviceTree_aw_bits_qos( outmemsys_io_deviceTree_aw_bits_qos ),
       .io_deviceTree_aw_bits_region( outmemsys_io_deviceTree_aw_bits_region ),
       .io_deviceTree_aw_bits_id( outmemsys_io_deviceTree_aw_bits_id ),
       .io_deviceTree_aw_bits_user( outmemsys_io_deviceTree_aw_bits_user ),
       .io_deviceTree_w_ready( deviceTree_io_w_ready ),
       .io_deviceTree_w_valid( outmemsys_io_deviceTree_w_valid ),
       .io_deviceTree_w_bits_data( outmemsys_io_deviceTree_w_bits_data ),
       .io_deviceTree_w_bits_last( outmemsys_io_deviceTree_w_bits_last ),
       .io_deviceTree_w_bits_strb( outmemsys_io_deviceTree_w_bits_strb ),
       .io_deviceTree_w_bits_user( outmemsys_io_deviceTree_w_bits_user ),
       .io_deviceTree_b_ready( outmemsys_io_deviceTree_b_ready ),
       .io_deviceTree_b_valid( deviceTree_io_b_valid ),
       //.io_deviceTree_b_bits_resp(  )
       //.io_deviceTree_b_bits_id(  )
       //.io_deviceTree_b_bits_user(  )
       .io_deviceTree_ar_ready( deviceTree_io_ar_ready ),
       .io_deviceTree_ar_valid( outmemsys_io_deviceTree_ar_valid ),
       .io_deviceTree_ar_bits_addr( outmemsys_io_deviceTree_ar_bits_addr ),
       .io_deviceTree_ar_bits_len( outmemsys_io_deviceTree_ar_bits_len ),
       .io_deviceTree_ar_bits_size( outmemsys_io_deviceTree_ar_bits_size ),
       .io_deviceTree_ar_bits_burst( outmemsys_io_deviceTree_ar_bits_burst ),
       .io_deviceTree_ar_bits_lock( outmemsys_io_deviceTree_ar_bits_lock ),
       .io_deviceTree_ar_bits_cache( outmemsys_io_deviceTree_ar_bits_cache ),
       .io_deviceTree_ar_bits_prot( outmemsys_io_deviceTree_ar_bits_prot ),
       .io_deviceTree_ar_bits_qos( outmemsys_io_deviceTree_ar_bits_qos ),
       .io_deviceTree_ar_bits_region( outmemsys_io_deviceTree_ar_bits_region ),
       .io_deviceTree_ar_bits_id( outmemsys_io_deviceTree_ar_bits_id ),
       .io_deviceTree_ar_bits_user( outmemsys_io_deviceTree_ar_bits_user ),
       .io_deviceTree_r_ready( outmemsys_io_deviceTree_r_ready ),
       .io_deviceTree_r_valid( deviceTree_io_r_valid ),
       .io_deviceTree_r_bits_resp( deviceTree_io_r_bits_resp ),
       .io_deviceTree_r_bits_data( deviceTree_io_r_bits_data ),
       .io_deviceTree_r_bits_last( deviceTree_io_r_bits_last ),
       .io_deviceTree_r_bits_id( deviceTree_io_r_bits_id ),
       .io_deviceTree_r_bits_user( deviceTree_io_r_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign outmemsys.io_mem_backup_req_bits = {1{$random}};
    assign outmemsys.io_deviceTree_b_bits_resp = {1{$random}};
    assign outmemsys.io_deviceTree_b_bits_id = {1{$random}};
    assign outmemsys.io_deviceTree_b_bits_user = {1{$random}};
// synthesis translate_on
`endif
  SmiArbiter_0 SmiArbiter(.clk(clk), .reset(reset),
       .io_in_1_req_ready( SmiArbiter_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_in_1_resp_valid( SmiArbiter_io_in_1_resp_valid ),
       .io_in_1_resp_bits( SmiArbiter_io_in_1_resp_bits ),
       .io_in_0_req_ready( SmiArbiter_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_in_0_resp_valid( SmiArbiter_io_in_0_resp_valid ),
       .io_in_0_resp_bits( SmiArbiter_io_in_0_resp_bits ),
       .io_out_req_ready( io_htif_0_csr_req_ready ),
       .io_out_req_valid( SmiArbiter_io_out_req_valid ),
       .io_out_req_bits_rw( SmiArbiter_io_out_req_bits_rw ),
       .io_out_req_bits_addr( SmiArbiter_io_out_req_bits_addr ),
       .io_out_req_bits_data( SmiArbiter_io_out_req_bits_data ),
       .io_out_resp_ready( SmiArbiter_io_out_resp_ready ),
       .io_out_resp_valid( io_htif_0_csr_resp_valid ),
       .io_out_resp_bits( io_htif_0_csr_resp_bits )
  );
  SCRFile scrFile(.clk(clk), .reset(reset),
       .io_smi_req_ready( scrFile_io_smi_req_ready ),
       .io_smi_req_valid( scrArb_io_out_req_valid ),
       .io_smi_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_smi_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_smi_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_smi_resp_ready( scrArb_io_out_resp_ready ),
       .io_smi_resp_valid( scrFile_io_smi_resp_valid ),
       .io_smi_resp_bits( scrFile_io_smi_resp_bits ),
       .io_scr_rdata_63( T34 ),
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       .io_scr_rdata_2( T12 ),
       .io_scr_rdata_1( 64'h400 ),
       .io_scr_rdata_0( 64'h1 ),
       .io_scr_wen( scrFile_io_scr_wen ),
       .io_scr_waddr( scrFile_io_scr_waddr ),
       .io_scr_wdata( scrFile_io_scr_wdata )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign scrFile.io_scr_rdata_62 = {2{$random}};
    assign scrFile.io_scr_rdata_61 = {2{$random}};
    assign scrFile.io_scr_rdata_60 = {2{$random}};
    assign scrFile.io_scr_rdata_59 = {2{$random}};
    assign scrFile.io_scr_rdata_58 = {2{$random}};
    assign scrFile.io_scr_rdata_57 = {2{$random}};
    assign scrFile.io_scr_rdata_56 = {2{$random}};
    assign scrFile.io_scr_rdata_55 = {2{$random}};
    assign scrFile.io_scr_rdata_54 = {2{$random}};
    assign scrFile.io_scr_rdata_53 = {2{$random}};
    assign scrFile.io_scr_rdata_52 = {2{$random}};
    assign scrFile.io_scr_rdata_51 = {2{$random}};
    assign scrFile.io_scr_rdata_50 = {2{$random}};
    assign scrFile.io_scr_rdata_49 = {2{$random}};
    assign scrFile.io_scr_rdata_48 = {2{$random}};
    assign scrFile.io_scr_rdata_47 = {2{$random}};
    assign scrFile.io_scr_rdata_46 = {2{$random}};
    assign scrFile.io_scr_rdata_45 = {2{$random}};
    assign scrFile.io_scr_rdata_44 = {2{$random}};
    assign scrFile.io_scr_rdata_43 = {2{$random}};
    assign scrFile.io_scr_rdata_42 = {2{$random}};
    assign scrFile.io_scr_rdata_41 = {2{$random}};
    assign scrFile.io_scr_rdata_40 = {2{$random}};
    assign scrFile.io_scr_rdata_39 = {2{$random}};
    assign scrFile.io_scr_rdata_38 = {2{$random}};
    assign scrFile.io_scr_rdata_37 = {2{$random}};
    assign scrFile.io_scr_rdata_36 = {2{$random}};
    assign scrFile.io_scr_rdata_35 = {2{$random}};
    assign scrFile.io_scr_rdata_34 = {2{$random}};
    assign scrFile.io_scr_rdata_33 = {2{$random}};
    assign scrFile.io_scr_rdata_32 = {2{$random}};
    assign scrFile.io_scr_rdata_31 = {2{$random}};
    assign scrFile.io_scr_rdata_30 = {2{$random}};
    assign scrFile.io_scr_rdata_29 = {2{$random}};
    assign scrFile.io_scr_rdata_28 = {2{$random}};
    assign scrFile.io_scr_rdata_27 = {2{$random}};
    assign scrFile.io_scr_rdata_26 = {2{$random}};
    assign scrFile.io_scr_rdata_25 = {2{$random}};
    assign scrFile.io_scr_rdata_24 = {2{$random}};
    assign scrFile.io_scr_rdata_23 = {2{$random}};
    assign scrFile.io_scr_rdata_22 = {2{$random}};
    assign scrFile.io_scr_rdata_21 = {2{$random}};
    assign scrFile.io_scr_rdata_20 = {2{$random}};
    assign scrFile.io_scr_rdata_19 = {2{$random}};
    assign scrFile.io_scr_rdata_18 = {2{$random}};
    assign scrFile.io_scr_rdata_17 = {2{$random}};
    assign scrFile.io_scr_rdata_16 = {2{$random}};
    assign scrFile.io_scr_rdata_15 = {2{$random}};
    assign scrFile.io_scr_rdata_14 = {2{$random}};
    assign scrFile.io_scr_rdata_13 = {2{$random}};
    assign scrFile.io_scr_rdata_12 = {2{$random}};
    assign scrFile.io_scr_rdata_11 = {2{$random}};
    assign scrFile.io_scr_rdata_10 = {2{$random}};
    assign scrFile.io_scr_rdata_9 = {2{$random}};
    assign scrFile.io_scr_rdata_8 = {2{$random}};
    assign scrFile.io_scr_rdata_7 = {2{$random}};
    assign scrFile.io_scr_rdata_6 = {2{$random}};
    assign scrFile.io_scr_rdata_5 = {2{$random}};
    assign scrFile.io_scr_rdata_4 = {2{$random}};
    assign scrFile.io_scr_rdata_3 = {2{$random}};
// synthesis translate_on
`endif
  SmiArbiter_1 scrArb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( scrArb_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_scr_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_in_1_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_in_0_req_ready( scrArb_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_scr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_scr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_scr_resp_ready ),
       .io_in_0_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( scrArb_io_in_0_resp_bits ),
       .io_out_req_ready( scrFile_io_smi_req_ready ),
       .io_out_req_valid( scrArb_io_out_req_valid ),
       .io_out_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_out_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_out_resp_ready( scrArb_io_out_resp_ready ),
       .io_out_resp_valid( scrFile_io_smi_resp_valid ),
       .io_out_resp_bits( scrFile_io_smi_resp_bits )
  );
  NastiROM deviceTree(.clk(clk), .reset(reset),
       .io_aw_ready( deviceTree_io_aw_ready ),
       .io_aw_valid( outmemsys_io_deviceTree_aw_valid ),
       .io_aw_bits_addr( outmemsys_io_deviceTree_aw_bits_addr ),
       .io_aw_bits_len( outmemsys_io_deviceTree_aw_bits_len ),
       .io_aw_bits_size( outmemsys_io_deviceTree_aw_bits_size ),
       .io_aw_bits_burst( outmemsys_io_deviceTree_aw_bits_burst ),
       .io_aw_bits_lock( outmemsys_io_deviceTree_aw_bits_lock ),
       .io_aw_bits_cache( outmemsys_io_deviceTree_aw_bits_cache ),
       .io_aw_bits_prot( outmemsys_io_deviceTree_aw_bits_prot ),
       .io_aw_bits_qos( outmemsys_io_deviceTree_aw_bits_qos ),
       .io_aw_bits_region( outmemsys_io_deviceTree_aw_bits_region ),
       .io_aw_bits_id( outmemsys_io_deviceTree_aw_bits_id ),
       .io_aw_bits_user( outmemsys_io_deviceTree_aw_bits_user ),
       .io_w_ready( deviceTree_io_w_ready ),
       .io_w_valid( outmemsys_io_deviceTree_w_valid ),
       .io_w_bits_data( outmemsys_io_deviceTree_w_bits_data ),
       .io_w_bits_last( outmemsys_io_deviceTree_w_bits_last ),
       .io_w_bits_strb( outmemsys_io_deviceTree_w_bits_strb ),
       .io_w_bits_user( outmemsys_io_deviceTree_w_bits_user ),
       .io_b_ready( outmemsys_io_deviceTree_b_ready ),
       .io_b_valid( deviceTree_io_b_valid ),
       //.io_b_bits_resp(  )
       //.io_b_bits_id(  )
       //.io_b_bits_user(  )
       .io_ar_ready( deviceTree_io_ar_ready ),
       .io_ar_valid( outmemsys_io_deviceTree_ar_valid ),
       .io_ar_bits_addr( outmemsys_io_deviceTree_ar_bits_addr ),
       .io_ar_bits_len( outmemsys_io_deviceTree_ar_bits_len ),
       .io_ar_bits_size( outmemsys_io_deviceTree_ar_bits_size ),
       .io_ar_bits_burst( outmemsys_io_deviceTree_ar_bits_burst ),
       .io_ar_bits_lock( outmemsys_io_deviceTree_ar_bits_lock ),
       .io_ar_bits_cache( outmemsys_io_deviceTree_ar_bits_cache ),
       .io_ar_bits_prot( outmemsys_io_deviceTree_ar_bits_prot ),
       .io_ar_bits_qos( outmemsys_io_deviceTree_ar_bits_qos ),
       .io_ar_bits_region( outmemsys_io_deviceTree_ar_bits_region ),
       .io_ar_bits_id( outmemsys_io_deviceTree_ar_bits_id ),
       .io_ar_bits_user( outmemsys_io_deviceTree_ar_bits_user ),
       .io_r_ready( outmemsys_io_deviceTree_r_ready ),
       .io_r_valid( deviceTree_io_r_valid ),
       .io_r_bits_resp( deviceTree_io_r_bits_resp ),
       .io_r_bits_data( deviceTree_io_r_bits_data ),
       .io_r_bits_last( deviceTree_io_r_bits_last ),
       .io_r_bits_id( deviceTree_io_r_bits_id ),
       .io_r_bits_user( deviceTree_io_r_bits_user )
  );
  SlowIO SlowIO(.clk(clk), .reset(reset),
       .io_out_fast_ready( SlowIO_io_out_fast_ready ),
       .io_out_fast_valid( T11 ),
       .io_out_fast_bits( T9 ),
       .io_out_slow_ready( T7 ),
       .io_out_slow_valid( SlowIO_io_out_slow_valid ),
       .io_out_slow_bits( SlowIO_io_out_slow_bits ),
       .io_in_fast_ready( T5 ),
       .io_in_fast_valid( SlowIO_io_in_fast_valid ),
       .io_in_fast_bits( SlowIO_io_in_fast_bits ),
       .io_in_slow_ready( SlowIO_io_in_slow_ready ),
       .io_in_slow_valid( T4 ),
       .io_in_slow_bits( T2 ),
       .io_clk_slow( SlowIO_io_clk_slow ),
       .io_set_divisor_valid( T0 ),
       .io_set_divisor_bits( T33 ),
       .io_divisor( SlowIO_io_divisor )
  );

  always @(posedge clk) begin
    if(T15) begin
      memory_channel_mux_select <= T14;
    end
    R29 <= T30;
    R32 <= io_host_clk;
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    input [11:0] io_rw_addr,
    input [2:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output io_csr_stall,
    output io_csr_xcpt,
    output io_eret,
    output io_status_sd,
    output[30:0] io_status_zero2,
    output io_status_sd_rv32,
    output[8:0] io_status_zero1,
    output[4:0] io_status_vm,
    output io_status_mprv,
    output[1:0] io_status_xs,
    output[1:0] io_status_fs,
    output[1:0] io_status_prv3,
    output io_status_ie3,
    output[1:0] io_status_prv2,
    output io_status_ie2,
    output[1:0] io_status_prv1,
    output io_status_ie1,
    output[1:0] io_status_prv,
    output io_status_ie,
    output[31:0] io_ptbr,
    output[39:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input [39:0] io_pc,
    output io_fatc,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [9:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[9:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[9:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_autl_acquire_ready
    input  io_rocc_autl_acquire_valid,
    input [25:0] io_rocc_autl_acquire_bits_addr_block,
    input [5:0] io_rocc_autl_acquire_bits_client_xact_id,
    input [1:0] io_rocc_autl_acquire_bits_addr_beat,
    input  io_rocc_autl_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_autl_acquire_bits_a_type,
    input [16:0] io_rocc_autl_acquire_bits_union,
    input [127:0] io_rocc_autl_acquire_bits_data,
    input  io_rocc_autl_grant_ready,
    //output io_rocc_autl_grant_valid
    //output[1:0] io_rocc_autl_grant_bits_addr_beat
    //output[5:0] io_rocc_autl_grant_bits_client_xact_id
    //output[3:0] io_rocc_autl_grant_bits_manager_xact_id
    //output io_rocc_autl_grant_bits_is_builtin_type
    //output[3:0] io_rocc_autl_grant_bits_g_type
    //output[127:0] io_rocc_autl_grant_bits_data
    //output io_rocc_fpu_req_ready
    input  io_rocc_fpu_req_valid,
    input [4:0] io_rocc_fpu_req_bits_cmd,
    input  io_rocc_fpu_req_bits_ldst,
    input  io_rocc_fpu_req_bits_wen,
    input  io_rocc_fpu_req_bits_ren1,
    input  io_rocc_fpu_req_bits_ren2,
    input  io_rocc_fpu_req_bits_ren3,
    input  io_rocc_fpu_req_bits_swap12,
    input  io_rocc_fpu_req_bits_swap23,
    input  io_rocc_fpu_req_bits_single,
    input  io_rocc_fpu_req_bits_fromint,
    input  io_rocc_fpu_req_bits_toint,
    input  io_rocc_fpu_req_bits_fastpipe,
    input  io_rocc_fpu_req_bits_fma,
    input  io_rocc_fpu_req_bits_div,
    input  io_rocc_fpu_req_bits_sqrt,
    input  io_rocc_fpu_req_bits_round,
    input  io_rocc_fpu_req_bits_wflags,
    input [2:0] io_rocc_fpu_req_bits_rm,
    input [1:0] io_rocc_fpu_req_bits_typ,
    input [64:0] io_rocc_fpu_req_bits_in1,
    input [64:0] io_rocc_fpu_req_bits_in2,
    input [64:0] io_rocc_fpu_req_bits_in3,
    input  io_rocc_fpu_resp_ready,
    //output io_rocc_fpu_resp_valid
    //output[64:0] io_rocc_fpu_resp_bits_data
    //output[4:0] io_rocc_fpu_resp_bits_exc
    //output io_rocc_exception
    output[11:0] io_rocc_csr_waddr,
    output[63:0] io_rocc_csr_wdata,
    output io_rocc_csr_wen,
    //output io_rocc_host_id
    output io_interrupt,
    output[63:0] io_interrupt_cause
);

  reg  T0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire csr_xcpt;
  wire insn_break;
  wire system_insn;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire insn_call;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire priv_sufficient;
  reg [1:0] reg_mstatus_prv;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  reg [1:0] reg_mstatus_prv1;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  reg [1:0] reg_mstatus_prv2;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[63:0] wdata;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [63:0] host_csr_bits_data;
  wire[63:0] T38;
  wire[63:0] T39;
  wire T40;
  wire host_csr_req_fire;
  wire T41;
  wire cpu_ren;
  wire T42;
  wire T43;
  reg  host_csr_req_valid;
  wire T44;
  wire T45;
  wire[63:0] T46;
  wire T47;
  wire[63:0] T48;
  wire[63:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire[11:0] addr;
  reg [11:0] host_csr_bits_addr;
  wire[11:0] T60;
  wire wen;
  wire T61;
  reg  host_csr_bits_rw;
  wire T62;
  wire T63;
  wire T64;
  wire read_only;
  wire[1:0] T65;
  wire cpu_wen;
  wire T66;
  wire T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T909;
  wire T75;
  wire T76;
  wire T77;
  wire insn_ret;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire insn_redirect_trap;
  wire maybe_insn_redirect_trap;
  wire T86;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[1:0] csr_addr_priv;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire fp_csr;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire addr_valid;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[1:0] T910;
  wire[2:0] T911;
  wire[1:0] T215;
  wire[1:0] T216;
  wire[1:0] T912;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] T220;
  wire[63:0] T221;
  wire[63:0] T222;
  wire T223;
  wire T224;
  wire T225;
  reg  reg_mstatus_ie;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg  reg_mstatus_ie1;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  reg  reg_mstatus_ie2;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  reg  reg_mip_ssip;
  wire T913;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  reg  reg_mie_ssip;
  wire T914;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  reg  reg_mip_msip;
  wire T915;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  reg  reg_mie_msip;
  wire T916;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  reg  reg_mip_stip;
  wire T917;
  wire T279;
  wire T280;
  reg  reg_mie_stip;
  wire T918;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  reg  reg_mip_mtip;
  wire T919;
  wire T291;
  wire T292;
  wire T293;
  reg [63:0] read_time;
  wire[63:0] T294;
  wire T295;
  reg [63:0] reg_mtimecmp;
  wire[63:0] T296;
  wire T297;
  reg  reg_mie_mtip;
  wire T920;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  reg [63:0] reg_fromhost;
  wire[63:0] T921;
  wire[63:0] T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  reg [2:0] reg_frm;
  wire[2:0] T922;
  wire[63:0] T318;
  wire[63:0] T319;
  wire[63:0] T923;
  wire T320;
  wire[63:0] T924;
  wire[58:0] T321;
  wire T322;
  wire[63:0] T323;
  reg [5:0] R324;
  wire[5:0] T925;
  wire[5:0] T325;
  wire[6:0] T326;
  wire[6:0] T926;
  reg [57:0] R327;
  wire[57:0] T927;
  wire[57:0] T328;
  wire[57:0] T329;
  wire T330;
  wire insn_sfence_vm;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire[39:0] T928;
  wire[63:0] T338;
  wire[63:0] T929;
  wire[39:0] T339;
  wire[39:0] T340;
  reg [39:0] reg_sepc;
  wire[39:0] T930;
  wire[63:0] T341;
  wire[63:0] T931;
  wire[39:0] T342;
  wire[63:0] T343;
  wire[63:0] T344;
  wire[63:0] T345;
  wire T346;
  reg [39:0] reg_mepc;
  wire[39:0] T932;
  wire[63:0] T347;
  wire[63:0] T933;
  wire[39:0] T348;
  wire[39:0] T349;
  wire[39:0] T350;
  wire[39:0] T351;
  wire[63:0] T352;
  wire[63:0] T353;
  wire[63:0] T354;
  wire T355;
  wire T356;
  wire[39:0] T357;
  reg [38:0] reg_stvec;
  wire[38:0] T934;
  wire[63:0] T358;
  wire[63:0] T935;
  wire[63:0] T359;
  wire[63:0] T360;
  wire[63:0] T361;
  wire T362;
  wire T363;
  wire[63:0] T364;
  reg [63:0] reg_mtvec;
  wire[63:0] T936;
  wire[63:0] T365;
  wire[63:0] T366;
  wire T367;
  wire[63:0] T937;
  wire[7:0] T368;
  wire T369;
  reg [31:0] reg_sptbr;
  wire[31:0] T370;
  wire[31:0] T371;
  wire[19:0] T372;
  wire T373;
  reg  reg_mstatus_ie3;
  wire T374;
  reg [1:0] reg_mstatus_prv3;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[1:0] T938;
  wire T377;
  reg [1:0] reg_mstatus_fs;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire[1:0] T382;
  wire[1:0] T383;
  wire[1:0] T939;
  wire T384;
  reg [1:0] reg_mstatus_xs;
  wire[1:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire[1:0] T389;
  reg  reg_mstatus_mprv;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  reg [4:0] reg_mstatus_vm;
  wire[4:0] T396;
  wire[4:0] T397;
  wire[4:0] T398;
  wire T399;
  wire T400;
  wire[4:0] T401;
  wire T402;
  wire T403;
  reg [8:0] reg_mstatus_zero1;
  wire[8:0] T404;
  reg  reg_mstatus_sd_rv32;
  wire T405;
  reg [30:0] reg_mstatus_zero2;
  wire[30:0] T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  reg  reg_wfi;
  wire T940;
  wire T411;
  wire T412;
  wire insn_wfi;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire some_interrupt_pending;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire[63:0] T437;
  wire[63:0] T438;
  wire[63:0] T439;
  wire[24:0] T440;
  wire[24:0] T941;
  wire T441;
  wire[63:0] T442;
  wire[63:0] T443;
  wire[63:0] T444;
  wire[23:0] T445;
  wire[23:0] T942;
  wire T446;
  wire[63:0] T447;
  wire[63:0] T448;
  wire[63:0] T943;
  wire[31:0] T449;
  wire[63:0] T450;
  wire[63:0] T451;
  wire[63:0] T452;
  reg [39:0] reg_sbadaddr;
  wire[39:0] T453;
  reg [39:0] reg_mbadaddr;
  wire[39:0] T454;
  wire[39:0] T455;
  wire[39:0] T456;
  wire[39:0] T457;
  wire[38:0] T458;
  wire T459;
  wire T460;
  wire[24:0] T461;
  wire T462;
  wire T463;
  wire[38:0] T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire[39:0] T473;
  wire T474;
  wire[23:0] T475;
  wire[23:0] T944;
  wire T476;
  wire[63:0] T477;
  wire[63:0] T478;
  reg [63:0] reg_scause;
  wire[63:0] T479;
  reg [63:0] reg_mcause;
  wire[63:0] T480;
  wire[63:0] T481;
  wire[63:0] T482;
  wire[63:0] T483;
  wire[63:0] T484;
  wire T485;
  wire T486;
  wire[63:0] T945;
  wire[3:0] T487;
  wire[3:0] T946;
  wire T488;
  wire[63:0] T489;
  wire T490;
  wire[63:0] T491;
  wire[63:0] T492;
  reg [63:0] reg_sscratch;
  wire[63:0] T493;
  wire T494;
  wire[63:0] T495;
  wire[63:0] T947;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[3:0] T499;
  wire[1:0] T500;
  wire T501;
  wire T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire[3:0] T506;
  wire[1:0] T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire T511;
  wire T512;
  wire[63:0] T513;
  wire[63:0] T948;
  wire[7:0] T514;
  wire[7:0] T515;
  wire[7:0] T516;
  wire[3:0] T517;
  wire[1:0] T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire T522;
  wire T523;
  wire[3:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire[1:0] T528;
  wire T529;
  wire T530;
  wire[63:0] T531;
  wire[63:0] T532;
  wire[63:0] T533;
  wire[63:0] T534;
  wire[13:0] T535;
  wire[3:0] T536;
  wire[2:0] T537;
  wire T538;
  wire T539;
  wire[63:0] read_mstatus;
  wire[63:0] T540;
  wire[11:0] T541;
  wire[5:0] T542;
  wire[2:0] T543;
  wire[2:0] T544;
  wire[5:0] T545;
  wire[2:0] T546;
  wire[2:0] T547;
  wire[51:0] T548;
  wire[9:0] T549;
  wire[3:0] T550;
  wire[5:0] T551;
  wire[41:0] T552;
  wire[9:0] T553;
  wire[31:0] T554;
  wire[1:0] T555;
  wire T556;
  wire T557;
  wire[9:0] T558;
  wire[7:0] T559;
  wire T560;
  wire T561;
  wire[6:0] T562;
  wire[1:0] T563;
  wire[1:0] T564;
  wire[49:0] T565;
  wire[16:0] T566;
  wire[2:0] T567;
  wire[1:0] T568;
  wire[1:0] T569;
  wire T570;
  wire T571;
  wire[13:0] T572;
  wire[32:0] T573;
  wire[31:0] T574;
  wire T575;
  wire T576;
  wire[30:0] T577;
  wire T578;
  wire T579;
  wire[63:0] T580;
  wire[63:0] T581;
  wire[63:0] T582;
  reg [5:0] R583;
  wire[5:0] T949;
  wire[5:0] T584;
  wire[5:0] T585;
  wire[6:0] T586;
  wire[6:0] T950;
  wire T587;
  reg [57:0] R588;
  wire[57:0] T951;
  wire[57:0] T589;
  wire[57:0] T590;
  wire T591;
  wire T592;
  wire[63:0] T593;
  wire[63:0] T594;
  wire[63:0] T595;
  reg [5:0] R596;
  wire[5:0] T952;
  wire[5:0] T597;
  wire[5:0] T598;
  wire[6:0] T599;
  wire[6:0] T953;
  wire T600;
  reg [57:0] R601;
  wire[57:0] T954;
  wire[57:0] T602;
  wire[57:0] T603;
  wire T604;
  wire T605;
  wire[63:0] T606;
  wire[63:0] T607;
  wire[63:0] T608;
  reg [5:0] R609;
  wire[5:0] T955;
  wire[5:0] T610;
  wire[5:0] T611;
  wire[6:0] T612;
  wire[6:0] T956;
  wire T613;
  reg [57:0] R614;
  wire[57:0] T957;
  wire[57:0] T615;
  wire[57:0] T616;
  wire T617;
  wire T618;
  wire[63:0] T619;
  wire[63:0] T620;
  wire[63:0] T621;
  reg [5:0] R622;
  wire[5:0] T958;
  wire[5:0] T623;
  wire[5:0] T624;
  wire[6:0] T625;
  wire[6:0] T959;
  wire T626;
  reg [57:0] R627;
  wire[57:0] T960;
  wire[57:0] T628;
  wire[57:0] T629;
  wire T630;
  wire T631;
  wire[63:0] T632;
  wire[63:0] T633;
  wire[63:0] T634;
  reg [5:0] R635;
  wire[5:0] T961;
  wire[5:0] T636;
  wire[5:0] T637;
  wire[6:0] T638;
  wire[6:0] T962;
  wire T639;
  reg [57:0] R640;
  wire[57:0] T963;
  wire[57:0] T641;
  wire[57:0] T642;
  wire T643;
  wire T644;
  wire[63:0] T645;
  wire[63:0] T646;
  wire[63:0] T647;
  reg [5:0] R648;
  wire[5:0] T964;
  wire[5:0] T649;
  wire[5:0] T650;
  wire[6:0] T651;
  wire[6:0] T965;
  wire T652;
  reg [57:0] R653;
  wire[57:0] T966;
  wire[57:0] T654;
  wire[57:0] T655;
  wire T656;
  wire T657;
  wire[63:0] T658;
  wire[63:0] T659;
  wire[63:0] T660;
  reg [5:0] R661;
  wire[5:0] T967;
  wire[5:0] T662;
  wire[5:0] T663;
  wire[6:0] T664;
  wire[6:0] T968;
  wire T665;
  reg [57:0] R666;
  wire[57:0] T969;
  wire[57:0] T667;
  wire[57:0] T668;
  wire T669;
  wire T670;
  wire[63:0] T671;
  wire[63:0] T672;
  wire[63:0] T673;
  reg [5:0] R674;
  wire[5:0] T970;
  wire[5:0] T675;
  wire[5:0] T676;
  wire[6:0] T677;
  wire[6:0] T971;
  wire T678;
  reg [57:0] R679;
  wire[57:0] T972;
  wire[57:0] T680;
  wire[57:0] T681;
  wire T682;
  wire T683;
  wire[63:0] T684;
  wire[63:0] T685;
  wire[63:0] T686;
  reg [5:0] R687;
  wire[5:0] T973;
  wire[5:0] T688;
  wire[5:0] T689;
  wire[6:0] T690;
  wire[6:0] T974;
  wire T691;
  reg [57:0] R692;
  wire[57:0] T975;
  wire[57:0] T693;
  wire[57:0] T694;
  wire T695;
  wire T696;
  wire[63:0] T697;
  wire[63:0] T698;
  wire[63:0] T699;
  reg [5:0] R700;
  wire[5:0] T976;
  wire[5:0] T701;
  wire[5:0] T702;
  wire[6:0] T703;
  wire[6:0] T977;
  wire T704;
  reg [57:0] R705;
  wire[57:0] T978;
  wire[57:0] T706;
  wire[57:0] T707;
  wire T708;
  wire T709;
  wire[63:0] T710;
  wire[63:0] T711;
  wire[63:0] T712;
  reg [5:0] R713;
  wire[5:0] T979;
  wire[5:0] T714;
  wire[5:0] T715;
  wire[6:0] T716;
  wire[6:0] T980;
  wire T717;
  reg [57:0] R718;
  wire[57:0] T981;
  wire[57:0] T719;
  wire[57:0] T720;
  wire T721;
  wire T722;
  wire[63:0] T723;
  wire[63:0] T724;
  wire[63:0] T725;
  reg [5:0] R726;
  wire[5:0] T982;
  wire[5:0] T727;
  wire[5:0] T728;
  wire[6:0] T729;
  wire[6:0] T983;
  wire T730;
  reg [57:0] R731;
  wire[57:0] T984;
  wire[57:0] T732;
  wire[57:0] T733;
  wire T734;
  wire T735;
  wire[63:0] T736;
  wire[63:0] T737;
  wire[63:0] T738;
  reg [5:0] R739;
  wire[5:0] T985;
  wire[5:0] T740;
  wire[5:0] T741;
  wire[6:0] T742;
  wire[6:0] T986;
  wire T743;
  reg [57:0] R744;
  wire[57:0] T987;
  wire[57:0] T745;
  wire[57:0] T746;
  wire T747;
  wire T748;
  wire[63:0] T749;
  wire[63:0] T750;
  wire[63:0] T751;
  reg [5:0] R752;
  wire[5:0] T988;
  wire[5:0] T753;
  wire[5:0] T754;
  wire[6:0] T755;
  wire[6:0] T989;
  wire T756;
  reg [57:0] R757;
  wire[57:0] T990;
  wire[57:0] T758;
  wire[57:0] T759;
  wire T760;
  wire T761;
  wire[63:0] T762;
  wire[63:0] T763;
  wire[63:0] T764;
  reg [5:0] R765;
  wire[5:0] T991;
  wire[5:0] T766;
  wire[5:0] T767;
  wire[6:0] T768;
  wire[6:0] T992;
  wire T769;
  reg [57:0] R770;
  wire[57:0] T993;
  wire[57:0] T771;
  wire[57:0] T772;
  wire T773;
  wire T774;
  wire[63:0] T775;
  wire[63:0] T776;
  wire[63:0] T777;
  reg [5:0] R778;
  wire[5:0] T994;
  wire[5:0] T779;
  wire[5:0] T780;
  wire[6:0] T781;
  wire[6:0] T995;
  wire T782;
  reg [57:0] R783;
  wire[57:0] T996;
  wire[57:0] T784;
  wire[57:0] T785;
  wire T786;
  wire T787;
  wire[63:0] T788;
  wire[63:0] T789;
  wire[63:0] T790;
  reg [5:0] R791;
  wire[5:0] T997;
  wire[5:0] T792;
  wire[5:0] T793;
  wire[5:0] T794;
  wire[6:0] T795;
  wire[6:0] T998;
  wire T796;
  wire[5:0] T797;
  wire T798;
  reg [57:0] R799;
  wire[57:0] T999;
  wire[57:0] T800;
  wire[57:0] T801;
  wire[57:0] T802;
  wire T803;
  wire T804;
  wire[57:0] T805;
  wire[63:0] T806;
  wire[63:0] T807;
  wire[63:0] T808;
  wire[63:0] T809;
  wire[63:0] T810;
  wire[63:0] T811;
  reg [63:0] reg_tohost;
  wire[63:0] T1000;
  wire[63:0] T812;
  wire[63:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire[63:0] T821;
  wire[63:0] T1001;
  wire T822;
  reg  reg_stats;
  wire T1002;
  wire T823;
  wire T824;
  wire T825;
  wire[63:0] T826;
  wire[63:0] T1003;
  wire T827;
  wire[63:0] T828;
  wire[63:0] T829;
  wire[63:0] T830;
  wire[63:0] T831;
  wire[63:0] T832;
  wire[63:0] T833;
  wire[63:0] T834;
  wire[23:0] T835;
  wire[23:0] T1004;
  wire T836;
  wire[63:0] T837;
  wire[63:0] T838;
  wire[63:0] T839;
  wire[23:0] T840;
  wire[23:0] T1005;
  wire T841;
  wire[63:0] T842;
  wire[63:0] T843;
  reg [63:0] reg_mscratch;
  wire[63:0] T844;
  wire T845;
  wire[63:0] T846;
  wire[63:0] T1006;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[3:0] T850;
  wire[1:0] T851;
  reg  reg_mie_usip;
  wire T1007;
  wire[1:0] T852;
  reg  reg_mie_hsip;
  wire T1008;
  wire[3:0] T853;
  wire[1:0] T854;
  reg  reg_mie_utip;
  wire T1009;
  wire[1:0] T855;
  reg  reg_mie_htip;
  wire T1010;
  wire[63:0] T856;
  wire[63:0] T1011;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[3:0] T860;
  wire[1:0] T861;
  reg  reg_mip_usip;
  wire T1012;
  wire[1:0] T862;
  reg  reg_mip_hsip;
  wire T1013;
  wire[3:0] T863;
  wire[1:0] T864;
  reg  reg_mip_utip;
  wire T1014;
  wire[1:0] T865;
  reg  reg_mip_htip;
  wire T1015;
  wire[63:0] T866;
  wire[63:0] T867;
  wire[63:0] T1016;
  wire[30:0] T868;
  wire[63:0] T869;
  wire[63:0] T870;
  wire[63:0] T871;
  wire[63:0] T872;
  wire[63:0] T873;
  wire[63:0] T874;
  wire[63:0] T875;
  wire[63:0] T1017;
  wire[63:0] T876;
  wire[63:0] T877;
  wire[63:0] T878;
  wire[63:0] T879;
  wire[63:0] T880;
  wire[63:0] T881;
  wire[63:0] T882;
  wire[63:0] T883;
  wire[63:0] T884;
  wire[63:0] T885;
  wire[63:0] T886;
  wire[63:0] T887;
  wire[63:0] T888;
  wire[63:0] T889;
  wire[63:0] T890;
  wire[63:0] T891;
  wire[63:0] T1018;
  wire[7:0] T892;
  wire[7:0] T893;
  wire[7:0] T894;
  reg [4:0] reg_fflags;
  wire[4:0] T1019;
  wire[63:0] T895;
  wire[63:0] T896;
  wire[63:0] T1020;
  wire[4:0] T897;
  wire[4:0] T898;
  wire T899;
  wire[7:0] T1021;
  wire[4:0] T900;
  wire[4:0] T1022;
  wire[2:0] T901;
  wire[4:0] T902;
  reg  host_csr_rep_valid;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    reg_mstatus_prv = {1{$random}};
    reg_mstatus_prv1 = {1{$random}};
    reg_mstatus_prv2 = {1{$random}};
    host_csr_bits_data = {2{$random}};
    host_csr_req_valid = {1{$random}};
    host_csr_bits_addr = {1{$random}};
    host_csr_bits_rw = {1{$random}};
    reg_mstatus_ie = {1{$random}};
    reg_mstatus_ie1 = {1{$random}};
    reg_mstatus_ie2 = {1{$random}};
    reg_mip_ssip = {1{$random}};
    reg_mie_ssip = {1{$random}};
    reg_mip_msip = {1{$random}};
    reg_mie_msip = {1{$random}};
    reg_mip_stip = {1{$random}};
    reg_mie_stip = {1{$random}};
    reg_mip_mtip = {1{$random}};
    read_time = {2{$random}};
    reg_mtimecmp = {2{$random}};
    reg_mie_mtip = {1{$random}};
    reg_fromhost = {2{$random}};
    reg_frm = {1{$random}};
    R324 = {1{$random}};
    R327 = {2{$random}};
    reg_sepc = {2{$random}};
    reg_mepc = {2{$random}};
    reg_stvec = {2{$random}};
    reg_mtvec = {2{$random}};
    reg_sptbr = {1{$random}};
    reg_mstatus_ie3 = {1{$random}};
    reg_mstatus_prv3 = {1{$random}};
    reg_mstatus_fs = {1{$random}};
    reg_mstatus_xs = {1{$random}};
    reg_mstatus_mprv = {1{$random}};
    reg_mstatus_vm = {1{$random}};
    reg_mstatus_zero1 = {1{$random}};
    reg_mstatus_sd_rv32 = {1{$random}};
    reg_mstatus_zero2 = {1{$random}};
    reg_wfi = {1{$random}};
    reg_sbadaddr = {2{$random}};
    reg_mbadaddr = {2{$random}};
    reg_scause = {2{$random}};
    reg_mcause = {2{$random}};
    reg_sscratch = {2{$random}};
    R583 = {1{$random}};
    R588 = {2{$random}};
    R596 = {1{$random}};
    R601 = {2{$random}};
    R609 = {1{$random}};
    R614 = {2{$random}};
    R622 = {1{$random}};
    R627 = {2{$random}};
    R635 = {1{$random}};
    R640 = {2{$random}};
    R648 = {1{$random}};
    R653 = {2{$random}};
    R661 = {1{$random}};
    R666 = {2{$random}};
    R674 = {1{$random}};
    R679 = {2{$random}};
    R687 = {1{$random}};
    R692 = {2{$random}};
    R700 = {1{$random}};
    R705 = {2{$random}};
    R713 = {1{$random}};
    R718 = {2{$random}};
    R726 = {1{$random}};
    R731 = {2{$random}};
    R739 = {1{$random}};
    R744 = {2{$random}};
    R752 = {1{$random}};
    R757 = {2{$random}};
    R765 = {1{$random}};
    R770 = {2{$random}};
    R778 = {1{$random}};
    R783 = {2{$random}};
    R791 = {1{$random}};
    R799 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_mscratch = {2{$random}};
    reg_mie_usip = {1{$random}};
    reg_mie_hsip = {1{$random}};
    reg_mie_utip = {1{$random}};
    reg_mie_htip = {1{$random}};
    reg_mip_usip = {1{$random}};
    reg_mip_hsip = {1{$random}};
    reg_mip_utip = {1{$random}};
    reg_mip_htip = {1{$random}};
    reg_fflags = {1{$random}};
    host_csr_rep_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_host_id = {1{$random}};
//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_fpu_resp_bits_exc = {1{$random}};
//  assign io_rocc_fpu_resp_bits_data = {3{$random}};
//  assign io_rocc_fpu_resp_valid = {1{$random}};
//  assign io_rocc_fpu_req_ready = {1{$random}};
//  assign io_rocc_autl_grant_bits_data = {4{$random}};
//  assign io_rocc_autl_grant_bits_g_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_autl_grant_valid = {1{$random}};
//  assign io_rocc_autl_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
//  assign io_rocc_cmd_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 <= 3'h1;
  assign T3 = T911 + T4;
  assign T4 = {1'h0, T5};
  assign T5 = T910 + T6;
  assign T6 = {1'h0, csr_xcpt};
  assign csr_xcpt = T11 | insn_break;
  assign insn_break = T7 & system_insn;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T7 = T9 & T8;
  assign T8 = io_rw_addr[1'h0];
  assign T9 = T10 ^ 1'h1;
  assign T10 = io_rw_addr[4'h8];
  assign T11 = T17 | insn_call;
  assign insn_call = T12 & system_insn;
  assign T12 = T15 & T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = io_rw_addr[1'h0];
  assign T15 = T16 ^ 1'h1;
  assign T16 = io_rw_addr[4'h8];
  assign T17 = T94 | T18;
  assign T18 = system_insn & T19;
  assign T19 = priv_sufficient ^ 1'h1;
  assign priv_sufficient = csr_addr_priv <= reg_mstatus_prv;
  assign T20 = reset ? 2'h3 : T21;
  assign T21 = T88 ? T87 : T22;
  assign T22 = insn_redirect_trap ? 2'h1 : T23;
  assign T23 = insn_ret ? reg_mstatus_prv1 : T24;
  assign T24 = T25 ? 2'h3 : reg_mstatus_prv;
  assign T25 = io_exception | csr_xcpt;
  assign T26 = reset ? 2'h3 : T27;
  assign T27 = T76 ? T909 : T28;
  assign T28 = T69 ? T68 : T29;
  assign T29 = insn_ret ? reg_mstatus_prv2 : T30;
  assign T30 = T25 ? reg_mstatus_prv : reg_mstatus_prv1;
  assign T31 = reset ? 2'h0 : T32;
  assign T32 = T52 ? T35 : T33;
  assign T33 = insn_ret ? 2'h0 : T34;
  assign T34 = T25 ? reg_mstatus_prv1 : reg_mstatus_prv2;
  assign T35 = wdata[4'h8:3'h7];
  assign wdata = T51 ? io_rw_wdata : T36;
  assign T36 = T50 ? T48 : T37;
  assign T37 = T47 ? T46 : host_csr_bits_data;
  assign T38 = host_csr_req_fire ? io_rw_rdata : T39;
  assign T39 = T40 ? io_host_csr_req_bits_data : host_csr_bits_data;
  assign T40 = io_host_csr_req_ready & io_host_csr_req_valid;
  assign host_csr_req_fire = host_csr_req_valid & T41;
  assign T41 = cpu_ren ^ 1'h1;
  assign cpu_ren = T43 & T42;
  assign T42 = system_insn ^ 1'h1;
  assign T43 = io_rw_cmd != 3'h0;
  assign T44 = host_csr_req_fire ? 1'h0 : T45;
  assign T45 = T40 ? 1'h1 : host_csr_req_valid;
  assign T46 = io_rw_rdata | io_rw_wdata;
  assign T47 = io_rw_cmd == 3'h2;
  assign T48 = io_rw_rdata & T49;
  assign T49 = ~ io_rw_wdata;
  assign T50 = io_rw_cmd == 3'h3;
  assign T51 = io_rw_cmd == 3'h1;
  assign T52 = T58 & T53;
  assign T53 = T55 | T54;
  assign T54 = 2'h1 == T35;
  assign T55 = T57 | T56;
  assign T56 = 2'h0 == T35;
  assign T57 = 2'h3 == T35;
  assign T58 = wen & T59;
  assign T59 = addr == 12'h300;
  assign addr = cpu_ren ? io_rw_addr : host_csr_bits_addr;
  assign T60 = T40 ? io_host_csr_req_bits_addr : host_csr_bits_addr;
  assign wen = T63 | T61;
  assign T61 = host_csr_req_fire & host_csr_bits_rw;
  assign T62 = T40 ? io_host_csr_req_bits_rw : host_csr_bits_rw;
  assign T63 = cpu_wen & T64;
  assign T64 = read_only ^ 1'h1;
  assign read_only = T65 == 2'h3;
  assign T65 = io_rw_addr[4'hb:4'ha];
  assign cpu_wen = T66 & priv_sufficient;
  assign T66 = cpu_ren & T67;
  assign T67 = io_rw_cmd != 3'h5;
  assign T68 = wdata[3'h5:3'h4];
  assign T69 = T58 & T70;
  assign T70 = T72 | T71;
  assign T71 = 2'h1 == T68;
  assign T72 = T74 | T73;
  assign T73 = 2'h0 == T68;
  assign T74 = 2'h3 == T68;
  assign T909 = {1'h0, T75};
  assign T75 = wdata[3'h4];
  assign T76 = wen & T77;
  assign T77 = addr == 12'h100;
  assign insn_ret = T78 & priv_sufficient;
  assign T78 = T79 & system_insn;
  assign T79 = T82 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_rw_addr[1'h0];
  assign T82 = T85 & T83;
  assign T83 = T84 ^ 1'h1;
  assign T84 = io_rw_addr[1'h1];
  assign T85 = io_rw_addr[4'h8];
  assign insn_redirect_trap = maybe_insn_redirect_trap & priv_sufficient;
  assign maybe_insn_redirect_trap = T86 & system_insn;
  assign T86 = io_rw_addr[2'h2];
  assign T87 = wdata[2'h2:1'h1];
  assign T88 = T58 & T89;
  assign T89 = T91 | T90;
  assign T90 = 2'h1 == T87;
  assign T91 = T93 | T92;
  assign T92 = 2'h0 == T87;
  assign T93 = 2'h3 == T87;
  assign csr_addr_priv = io_rw_addr[4'h9:4'h8];
  assign T94 = T214 | T95;
  assign T95 = cpu_ren & T96;
  assign T96 = T104 | T97;
  assign T97 = fp_csr & T98;
  assign T98 = T99 ^ 1'h1;
  assign T99 = io_status_fs != 2'h0;
  assign fp_csr = T101 | T100;
  assign T100 = addr == 12'h3;
  assign T101 = T103 | T102;
  assign T102 = addr == 12'h2;
  assign T103 = addr == 12'h1;
  assign T104 = T213 | T105;
  assign T105 = addr_valid ^ 1'h1;
  assign addr_valid = T107 | T106;
  assign T106 = addr == 12'h101;
  assign T107 = T109 | T108;
  assign T108 = addr == 12'h141;
  assign T109 = T111 | T110;
  assign T110 = addr == 12'h181;
  assign T111 = T113 | T112;
  assign T112 = addr == 12'h180;
  assign T113 = T115 | T114;
  assign T114 = addr == 12'hd43;
  assign T115 = T117 | T116;
  assign T116 = addr == 12'hd42;
  assign T117 = T119 | T118;
  assign T118 = addr == 12'h140;
  assign T119 = T121 | T120;
  assign T120 = addr == 12'h104;
  assign T121 = T123 | T122;
  assign T122 = addr == 12'h144;
  assign T123 = T124 | T77;
  assign T124 = T126 | T125;
  assign T125 = addr == 12'hccf;
  assign T126 = T128 | T127;
  assign T127 = addr == 12'hcce;
  assign T128 = T130 | T129;
  assign T129 = addr == 12'hccd;
  assign T130 = T132 | T131;
  assign T131 = addr == 12'hccc;
  assign T132 = T134 | T133;
  assign T133 = addr == 12'hccb;
  assign T134 = T136 | T135;
  assign T135 = addr == 12'hcca;
  assign T136 = T138 | T137;
  assign T137 = addr == 12'hcc9;
  assign T138 = T140 | T139;
  assign T139 = addr == 12'hcc8;
  assign T140 = T142 | T141;
  assign T141 = addr == 12'hcc7;
  assign T142 = T144 | T143;
  assign T143 = addr == 12'hcc6;
  assign T144 = T146 | T145;
  assign T145 = addr == 12'hcc5;
  assign T146 = T148 | T147;
  assign T147 = addr == 12'hcc4;
  assign T148 = T150 | T149;
  assign T149 = addr == 12'hcc3;
  assign T150 = T152 | T151;
  assign T151 = addr == 12'hcc2;
  assign T152 = T154 | T153;
  assign T153 = addr == 12'hcc1;
  assign T154 = T156 | T155;
  assign T155 = addr == 12'hcc0;
  assign T156 = T158 | T157;
  assign T157 = addr == 12'h902;
  assign T158 = T160 | T159;
  assign T159 = addr == 12'hc02;
  assign T160 = T162 | T161;
  assign T161 = addr == 12'h781;
  assign T162 = T164 | T163;
  assign T163 = addr == 12'h780;
  assign T164 = T166 | T165;
  assign T165 = addr == 12'hc0;
  assign T166 = T168 | T167;
  assign T167 = addr == 12'hf10;
  assign T168 = T170 | T169;
  assign T169 = addr == 12'h321;
  assign T170 = T172 | T171;
  assign T171 = addr == 12'h342;
  assign T172 = T174 | T173;
  assign T173 = addr == 12'h343;
  assign T174 = T176 | T175;
  assign T175 = addr == 12'h341;
  assign T176 = T178 | T177;
  assign T177 = addr == 12'h340;
  assign T178 = T180 | T179;
  assign T179 = addr == 12'h304;
  assign T180 = T182 | T181;
  assign T181 = addr == 12'h344;
  assign T182 = T184 | T183;
  assign T183 = addr == 12'h783;
  assign T184 = T186 | T185;
  assign T185 = addr == 12'h784;
  assign T186 = T188 | T187;
  assign T187 = addr == 12'h301;
  assign T188 = T190 | T189;
  assign T189 = addr == 12'h782;
  assign T190 = T192 | T191;
  assign T191 = addr == 12'h302;
  assign T192 = T193 | T59;
  assign T193 = T195 | T194;
  assign T194 = addr == 12'hf01;
  assign T195 = T197 | T196;
  assign T196 = addr == 12'hf00;
  assign T197 = T199 | T198;
  assign T198 = addr == 12'h701;
  assign T199 = T201 | T200;
  assign T200 = addr == 12'ha01;
  assign T201 = T203 | T202;
  assign T202 = addr == 12'hd01;
  assign T203 = T205 | T204;
  assign T204 = addr == 12'h901;
  assign T205 = T207 | T206;
  assign T206 = addr == 12'hc01;
  assign T207 = T209 | T208;
  assign T208 = addr == 12'h900;
  assign T209 = T211 | T210;
  assign T210 = addr == 12'hc00;
  assign T211 = T212 | T100;
  assign T212 = T103 | T102;
  assign T213 = priv_sufficient ^ 1'h1;
  assign T214 = cpu_wen & read_only;
  assign T910 = {1'h0, io_exception};
  assign T911 = {1'h0, T215};
  assign T215 = T912 + T216;
  assign T216 = {1'h0, insn_redirect_trap};
  assign T912 = {1'h0, insn_ret};
  assign io_interrupt_cause = T217;
  assign T217 = T312 ? 64'h8000000000000003 : T218;
  assign T218 = T300 ? 64'h8000000000000002 : T219;
  assign T219 = T285 ? 64'h8000000000000001 : T220;
  assign T220 = T273 ? 64'h8000000000000001 : T221;
  assign T221 = T260 ? 64'h8000000000000000 : T222;
  assign T222 = T223 ? 64'h8000000000000000 : 64'h0;
  assign T223 = T247 & T224;
  assign T224 = T246 | T225;
  assign T225 = T245 & reg_mstatus_ie;
  assign T226 = reset ? 1'h0 : T227;
  assign T227 = T76 ? T244 : T228;
  assign T228 = T58 ? T243 : T229;
  assign T229 = insn_ret ? reg_mstatus_ie1 : T230;
  assign T230 = T25 ? 1'h0 : reg_mstatus_ie;
  assign T231 = reset ? 1'h0 : T232;
  assign T232 = T76 ? T242 : T233;
  assign T233 = T58 ? T241 : T234;
  assign T234 = insn_ret ? reg_mstatus_ie2 : T235;
  assign T235 = T25 ? reg_mstatus_ie : reg_mstatus_ie1;
  assign T236 = reset ? 1'h0 : T237;
  assign T237 = T58 ? T240 : T238;
  assign T238 = insn_ret ? 1'h1 : T239;
  assign T239 = T25 ? reg_mstatus_ie1 : reg_mstatus_ie2;
  assign T240 = wdata[3'h6];
  assign T241 = wdata[2'h3];
  assign T242 = wdata[2'h3];
  assign T243 = wdata[1'h0];
  assign T244 = wdata[1'h0];
  assign T245 = reg_mstatus_prv == 2'h1;
  assign T246 = reg_mstatus_prv < 2'h1;
  assign T247 = reg_mie_ssip & reg_mip_ssip;
  assign T913 = reset ? 1'h0 : T248;
  assign T248 = T253 ? T252 : T249;
  assign T249 = T251 ? T250 : reg_mip_ssip;
  assign T250 = wdata[1'h1];
  assign T251 = wen & T181;
  assign T252 = wdata[1'h1];
  assign T253 = wen & T122;
  assign T914 = reset ? 1'h0 : T254;
  assign T254 = T259 ? T258 : T255;
  assign T255 = T257 ? T256 : reg_mie_ssip;
  assign T256 = wdata[1'h1];
  assign T257 = wen & T179;
  assign T258 = wdata[1'h1];
  assign T259 = wen & T120;
  assign T260 = T265 & T261;
  assign T261 = T264 | T262;
  assign T262 = T263 & reg_mstatus_ie;
  assign T263 = reg_mstatus_prv == 2'h3;
  assign T264 = reg_mstatus_prv < 2'h3;
  assign T265 = reg_mie_msip & reg_mip_msip;
  assign T915 = reset ? 1'h0 : T266;
  assign T266 = T270 ? T269 : T267;
  assign T267 = T251 ? T268 : reg_mip_msip;
  assign T268 = wdata[2'h3];
  assign T269 = wdata[1'h0];
  assign T270 = wen & T183;
  assign T916 = reset ? 1'h0 : T271;
  assign T271 = T257 ? T272 : reg_mie_msip;
  assign T272 = wdata[2'h3];
  assign T273 = T278 & T274;
  assign T274 = T277 | T275;
  assign T275 = T276 & reg_mstatus_ie;
  assign T276 = reg_mstatus_prv == 2'h1;
  assign T277 = reg_mstatus_prv < 2'h1;
  assign T278 = reg_mie_stip & reg_mip_stip;
  assign T917 = reset ? 1'h0 : T279;
  assign T279 = T251 ? T280 : reg_mip_stip;
  assign T280 = wdata[3'h5];
  assign T918 = reset ? 1'h0 : T281;
  assign T281 = T259 ? T284 : T282;
  assign T282 = T257 ? T283 : reg_mie_stip;
  assign T283 = wdata[3'h5];
  assign T284 = wdata[3'h5];
  assign T285 = T290 & T286;
  assign T286 = T289 | T287;
  assign T287 = T288 & reg_mstatus_ie;
  assign T288 = reg_mstatus_prv == 2'h3;
  assign T289 = reg_mstatus_prv < 2'h3;
  assign T290 = reg_mie_mtip & reg_mip_mtip;
  assign T919 = reset ? 1'h0 : T291;
  assign T291 = T297 ? 1'h0 : T292;
  assign T292 = T293 ? 1'h1 : reg_mip_mtip;
  assign T293 = reg_mtimecmp <= read_time;
  assign T294 = T295 ? wdata : read_time;
  assign T295 = wen & T198;
  assign T296 = T297 ? wdata : reg_mtimecmp;
  assign T297 = wen & T169;
  assign T920 = reset ? 1'h0 : T298;
  assign T298 = T257 ? T299 : reg_mie_mtip;
  assign T299 = wdata[3'h7];
  assign T300 = T305 & T301;
  assign T301 = T304 | T302;
  assign T302 = T303 & reg_mstatus_ie;
  assign T303 = reg_mstatus_prv == 2'h3;
  assign T304 = reg_mstatus_prv < 2'h3;
  assign T305 = reg_fromhost != 64'h0;
  assign T921 = reset ? 64'h0 : T306;
  assign T306 = T307 ? wdata : reg_fromhost;
  assign T307 = T311 & T308;
  assign T308 = T310 | T309;
  assign T309 = host_csr_req_fire ^ 1'h1;
  assign T310 = reg_fromhost == 64'h0;
  assign T311 = wen & T161;
  assign T312 = io_rocc_interrupt & T313;
  assign T313 = T316 | T314;
  assign T314 = T315 & reg_mstatus_ie;
  assign T315 = reg_mstatus_prv == 2'h3;
  assign T316 = reg_mstatus_prv < 2'h3;
  assign io_interrupt = T317;
  assign T317 = io_interrupt_cause[6'h3f];
  assign io_rocc_csr_wen = wen;
  assign io_rocc_csr_wdata = wdata;
  assign io_rocc_csr_waddr = addr;
  assign io_fcsr_rm = reg_frm;
  assign T922 = T318[2'h2:1'h0];
  assign T318 = T322 ? T924 : T319;
  assign T319 = T320 ? wdata : T923;
  assign T923 = {61'h0, reg_frm};
  assign T320 = wen & T102;
  assign T924 = {5'h0, T321};
  assign T321 = wdata >> 3'h5;
  assign T322 = wen & T100;
  assign io_time = T323;
  assign T323 = {R327, R324};
  assign T925 = reset ? 6'h0 : T325;
  assign T325 = T326[3'h5:1'h0];
  assign T326 = T926 + 7'h1;
  assign T926 = {1'h0, R324};
  assign T927 = reset ? 58'h0 : T328;
  assign T328 = T330 ? T329 : R327;
  assign T329 = R327 + 58'h1;
  assign T330 = T326[3'h6];
  assign io_fatc = insn_sfence_vm;
  assign insn_sfence_vm = T331 & priv_sufficient;
  assign T331 = T332 & system_insn;
  assign T332 = T334 & T333;
  assign T333 = io_rw_addr[1'h0];
  assign T334 = T337 & T335;
  assign T335 = T336 ^ 1'h1;
  assign T336 = io_rw_addr[1'h1];
  assign T337 = io_rw_addr[4'h8];
  assign io_evec = T928;
  assign T928 = T338[6'h27:1'h0];
  assign T338 = T369 ? T364 : T929;
  assign T929 = {24'h0, T339};
  assign T339 = maybe_insn_redirect_trap ? T357 : T340;
  assign T340 = T356 ? reg_mepc : reg_sepc;
  assign T930 = T341[6'h27:1'h0];
  assign T341 = T346 ? T343 : T931;
  assign T931 = {24'h0, T342};
  assign T342 = insn_redirect_trap ? reg_mepc : reg_sepc;
  assign T343 = ~ T344;
  assign T344 = T345 | 64'h3;
  assign T345 = ~ wdata;
  assign T346 = wen & T108;
  assign T932 = T347[6'h27:1'h0];
  assign T347 = T355 ? T352 : T933;
  assign T933 = {24'h0, T348};
  assign T348 = T25 ? T349 : reg_mepc;
  assign T349 = ~ T350;
  assign T350 = T351 | 40'h3;
  assign T351 = ~ io_pc;
  assign T352 = ~ T353;
  assign T353 = T354 | 64'h3;
  assign T354 = ~ wdata;
  assign T355 = wen & T175;
  assign T356 = reg_mstatus_prv[1'h1];
  assign T357 = {T363, reg_stvec};
  assign T934 = T358[6'h26:1'h0];
  assign T358 = T362 ? T359 : T935;
  assign T935 = {25'h0, reg_stvec};
  assign T359 = ~ T360;
  assign T360 = T361 | 64'h3;
  assign T361 = ~ wdata;
  assign T362 = wen & T106;
  assign T363 = reg_stvec[6'h26];
  assign T364 = T937 + reg_mtvec;
  assign T936 = reset ? 64'h100 : T365;
  assign T365 = T367 ? T366 : reg_mtvec;
  assign T366 = wdata & 64'h0;
  assign T367 = wen & T187;
  assign T937 = {56'h0, T368};
  assign T368 = reg_mstatus_prv << 3'h6;
  assign T369 = io_exception | csr_xcpt;
  assign io_ptbr = reg_sptbr;
  assign T370 = T373 ? T371 : reg_sptbr;
  assign T371 = {T372, 12'h0};
  assign T372 = wdata[5'h1f:4'hc];
  assign T373 = wen & T112;
  assign io_status_ie = reg_mstatus_ie;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_ie1 = reg_mstatus_ie1;
  assign io_status_prv1 = reg_mstatus_prv1;
  assign io_status_ie2 = reg_mstatus_ie2;
  assign io_status_prv2 = reg_mstatus_prv2;
  assign io_status_ie3 = reg_mstatus_ie3;
  assign T374 = reset ? 1'h0 : reg_mstatus_ie3;
  assign io_status_prv3 = reg_mstatus_prv3;
  assign T375 = reset ? 2'h0 : reg_mstatus_prv3;
  assign io_status_fs = T376;
  assign T376 = 2'h0 - T938;
  assign T938 = {1'h0, T377};
  assign T377 = reg_mstatus_fs != 2'h0;
  assign T378 = reset ? 2'h0 : T379;
  assign T379 = T76 ? T382 : T380;
  assign T380 = T58 ? T381 : reg_mstatus_fs;
  assign T381 = wdata[4'hd:4'hc];
  assign T382 = wdata[4'hd:4'hc];
  assign io_status_xs = T383;
  assign T383 = 2'h0 - T939;
  assign T939 = {1'h0, T384};
  assign T384 = reg_mstatus_xs != 2'h0;
  assign T385 = reset ? 2'h0 : T386;
  assign T386 = T76 ? T389 : T387;
  assign T387 = T58 ? T388 : reg_mstatus_xs;
  assign T388 = wdata[4'hf:4'he];
  assign T389 = wdata[4'hf:4'he];
  assign io_status_mprv = reg_mstatus_mprv;
  assign T390 = reset ? 1'h0 : T391;
  assign T391 = T76 ? T395 : T392;
  assign T392 = T58 ? T394 : T393;
  assign T393 = T25 ? 1'h0 : reg_mstatus_mprv;
  assign T394 = wdata[5'h10];
  assign T395 = wdata[5'h10];
  assign io_status_vm = reg_mstatus_vm;
  assign T396 = reset ? 5'h0 : T397;
  assign T397 = T402 ? 5'h9 : T398;
  assign T398 = T399 ? 5'h0 : reg_mstatus_vm;
  assign T399 = T58 & T400;
  assign T400 = T401 == 5'h0;
  assign T401 = wdata[5'h15:5'h11];
  assign T402 = T58 & T403;
  assign T403 = T401 == 5'h9;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign T404 = reset ? 9'h0 : reg_mstatus_zero1;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign T405 = reset ? 1'h0 : reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign T406 = reset ? 31'h0 : reg_mstatus_zero2;
  assign io_status_sd = T407;
  assign T407 = T409 | T408;
  assign T408 = io_status_xs == 2'h3;
  assign T409 = io_status_fs == 2'h3;
  assign io_eret = T410;
  assign T410 = insn_ret | insn_redirect_trap;
  assign io_csr_xcpt = csr_xcpt;
  assign io_csr_stall = reg_wfi;
  assign T940 = reset ? 1'h0 : T411;
  assign T411 = some_interrupt_pending ? 1'h0 : T412;
  assign T412 = insn_wfi ? 1'h1 : reg_wfi;
  assign insn_wfi = T413 & priv_sufficient;
  assign T413 = T414 & system_insn;
  assign T414 = T417 & T415;
  assign T415 = T416 ^ 1'h1;
  assign T416 = io_rw_addr[1'h0];
  assign T417 = T419 & T418;
  assign T418 = io_rw_addr[1'h1];
  assign T419 = io_rw_addr[4'h8];
  assign some_interrupt_pending = T420;
  assign T420 = T435 ? 1'h1 : T421;
  assign T421 = T433 ? 1'h1 : T422;
  assign T422 = T431 ? 1'h1 : T423;
  assign T423 = T429 ? 1'h1 : T424;
  assign T424 = T427 ? 1'h1 : T425;
  assign T425 = T247 & T426;
  assign T426 = reg_mstatus_prv <= 2'h1;
  assign T427 = T265 & T428;
  assign T428 = reg_mstatus_prv <= 2'h3;
  assign T429 = T278 & T430;
  assign T430 = reg_mstatus_prv <= 2'h1;
  assign T431 = T290 & T432;
  assign T432 = reg_mstatus_prv <= 2'h3;
  assign T433 = T305 & T434;
  assign T434 = reg_mstatus_prv <= 2'h3;
  assign T435 = io_rocc_interrupt & T436;
  assign T436 = reg_mstatus_prv <= 2'h3;
  assign io_rw_rdata = T437;
  assign T437 = T442 | T438;
  assign T438 = T106 ? T439 : 64'h0;
  assign T439 = {T440, reg_stvec};
  assign T440 = 25'h0 - T941;
  assign T941 = {24'h0, T441};
  assign T441 = reg_stvec[6'h26];
  assign T442 = T447 | T443;
  assign T443 = T108 ? T444 : 64'h0;
  assign T444 = {T445, reg_sepc};
  assign T445 = 24'h0 - T942;
  assign T942 = {23'h0, T446};
  assign T446 = reg_sepc[6'h27];
  assign T447 = T448 | 64'h0;
  assign T448 = T450 | T943;
  assign T943 = {32'h0, T449};
  assign T449 = T112 ? reg_sptbr : 32'h0;
  assign T450 = T477 | T451;
  assign T451 = T114 ? T452 : 64'h0;
  assign T452 = {T475, reg_sbadaddr};
  assign T453 = insn_redirect_trap ? reg_mbadaddr : reg_sbadaddr;
  assign T454 = T474 ? T473 : T455;
  assign T455 = T465 ? T457 : T456;
  assign T456 = T25 ? io_pc : reg_mbadaddr;
  assign T457 = {T459, T458};
  assign T458 = io_rw_wdata[6'h26:1'h0];
  assign T459 = T463 ? T462 : T460;
  assign T460 = T461 != 25'h0;
  assign T461 = io_rw_wdata[6'h3f:6'h27];
  assign T462 = T461 == 25'h1ffffff;
  assign T463 = $signed(T464) < $signed(1'h0);
  assign T464 = T458;
  assign T465 = T25 & T466;
  assign T466 = T468 | T467;
  assign T467 = io_cause == 64'h6;
  assign T468 = T470 | T469;
  assign T469 = io_cause == 64'h7;
  assign T470 = T472 | T471;
  assign T471 = io_cause == 64'h4;
  assign T472 = io_cause == 64'h5;
  assign T473 = wdata[6'h27:1'h0];
  assign T474 = wen & T173;
  assign T475 = 24'h0 - T944;
  assign T944 = {23'h0, T476};
  assign T476 = reg_sbadaddr[6'h27];
  assign T477 = T491 | T478;
  assign T478 = T116 ? reg_scause : 64'h0;
  assign T479 = insn_redirect_trap ? reg_mcause : reg_scause;
  assign T480 = T490 ? T489 : T481;
  assign T481 = T488 ? T945 : T482;
  assign T482 = T486 ? 64'h3 : T483;
  assign T483 = T485 ? 64'h2 : T484;
  assign T484 = T25 ? io_cause : reg_mcause;
  assign T485 = T25 & csr_xcpt;
  assign T486 = T485 & insn_break;
  assign T945 = {60'h0, T487};
  assign T487 = T946 + 4'h8;
  assign T946 = {2'h0, reg_mstatus_prv};
  assign T488 = T485 & insn_call;
  assign T489 = wdata & 64'h800000000000001f;
  assign T490 = wen & T171;
  assign T491 = T495 | T492;
  assign T492 = T118 ? reg_sscratch : 64'h0;
  assign T493 = T494 ? wdata : reg_sscratch;
  assign T494 = wen & T118;
  assign T495 = T513 | T947;
  assign T947 = {56'h0, T496};
  assign T496 = T120 ? T497 : 8'h0;
  assign T497 = T498;
  assign T498 = {T506, T499};
  assign T499 = {T503, T500};
  assign T500 = {T502, T501};
  assign T501 = 1'h0;
  assign T502 = reg_mie_ssip;
  assign T503 = {T505, T504};
  assign T504 = 1'h0;
  assign T505 = 1'h0;
  assign T506 = {T510, T507};
  assign T507 = {T509, T508};
  assign T508 = 1'h0;
  assign T509 = reg_mie_stip;
  assign T510 = {T512, T511};
  assign T511 = 1'h0;
  assign T512 = 1'h0;
  assign T513 = T531 | T948;
  assign T948 = {56'h0, T514};
  assign T514 = T122 ? T515 : 8'h0;
  assign T515 = T516;
  assign T516 = {T524, T517};
  assign T517 = {T521, T518};
  assign T518 = {T520, T519};
  assign T519 = 1'h0;
  assign T520 = reg_mip_ssip;
  assign T521 = {T523, T522};
  assign T522 = 1'h0;
  assign T523 = 1'h0;
  assign T524 = {T528, T525};
  assign T525 = {T527, T526};
  assign T526 = 1'h0;
  assign T527 = reg_mip_stip;
  assign T528 = {T530, T529};
  assign T529 = 1'h0;
  assign T530 = 1'h0;
  assign T531 = T580 | T532;
  assign T532 = T77 ? T533 : 64'h0;
  assign T533 = T534;
  assign T534 = {T565, T535};
  assign T535 = {T558, T536};
  assign T536 = {T556, T537};
  assign T537 = {T555, T538};
  assign T538 = T539;
  assign T539 = read_mstatus[1'h0];
  assign read_mstatus = T540;
  assign T540 = {T548, T541};
  assign T541 = {T545, T542};
  assign T542 = {T544, T543};
  assign T543 = {io_status_prv, io_status_ie};
  assign T544 = {io_status_prv1, io_status_ie1};
  assign T545 = {T547, T546};
  assign T546 = {io_status_prv2, io_status_ie2};
  assign T547 = {io_status_prv3, io_status_ie3};
  assign T548 = {T552, T549};
  assign T549 = {T551, T550};
  assign T550 = {io_status_xs, io_status_fs};
  assign T551 = {io_status_vm, io_status_mprv};
  assign T552 = {T554, T553};
  assign T553 = {io_status_sd_rv32, io_status_zero1};
  assign T554 = {io_status_sd, io_status_zero2};
  assign T555 = 2'h0;
  assign T556 = T557;
  assign T557 = read_mstatus[2'h3];
  assign T558 = {T563, T559};
  assign T559 = {T562, T560};
  assign T560 = T561;
  assign T561 = read_mstatus[3'h4];
  assign T562 = 7'h0;
  assign T563 = T564;
  assign T564 = read_mstatus[4'hd:4'hc];
  assign T565 = {T573, T566};
  assign T566 = {T572, T567};
  assign T567 = {T570, T568};
  assign T568 = T569;
  assign T569 = read_mstatus[4'hf:4'he];
  assign T570 = T571;
  assign T571 = read_mstatus[5'h10];
  assign T572 = 14'h0;
  assign T573 = {T578, T574};
  assign T574 = {T577, T575};
  assign T575 = T576;
  assign T576 = read_mstatus[5'h1f];
  assign T577 = 31'h0;
  assign T578 = T579;
  assign T579 = read_mstatus[6'h3f];
  assign T580 = T593 | T581;
  assign T581 = T125 ? T582 : 64'h0;
  assign T582 = {R588, R583};
  assign T949 = reset ? 6'h0 : T584;
  assign T584 = T587 ? T585 : R583;
  assign T585 = T586[3'h5:1'h0];
  assign T586 = T950 + 7'h1;
  assign T950 = {1'h0, R583};
  assign T587 = io_uarch_counters_15 != 1'h0;
  assign T951 = reset ? 58'h0 : T589;
  assign T589 = T591 ? T590 : R588;
  assign T590 = R588 + 58'h1;
  assign T591 = T587 & T592;
  assign T592 = T586[3'h6];
  assign T593 = T606 | T594;
  assign T594 = T127 ? T595 : 64'h0;
  assign T595 = {R601, R596};
  assign T952 = reset ? 6'h0 : T597;
  assign T597 = T600 ? T598 : R596;
  assign T598 = T599[3'h5:1'h0];
  assign T599 = T953 + 7'h1;
  assign T953 = {1'h0, R596};
  assign T600 = io_uarch_counters_14 != 1'h0;
  assign T954 = reset ? 58'h0 : T602;
  assign T602 = T604 ? T603 : R601;
  assign T603 = R601 + 58'h1;
  assign T604 = T600 & T605;
  assign T605 = T599[3'h6];
  assign T606 = T619 | T607;
  assign T607 = T129 ? T608 : 64'h0;
  assign T608 = {R614, R609};
  assign T955 = reset ? 6'h0 : T610;
  assign T610 = T613 ? T611 : R609;
  assign T611 = T612[3'h5:1'h0];
  assign T612 = T956 + 7'h1;
  assign T956 = {1'h0, R609};
  assign T613 = io_uarch_counters_13 != 1'h0;
  assign T957 = reset ? 58'h0 : T615;
  assign T615 = T617 ? T616 : R614;
  assign T616 = R614 + 58'h1;
  assign T617 = T613 & T618;
  assign T618 = T612[3'h6];
  assign T619 = T632 | T620;
  assign T620 = T131 ? T621 : 64'h0;
  assign T621 = {R627, R622};
  assign T958 = reset ? 6'h0 : T623;
  assign T623 = T626 ? T624 : R622;
  assign T624 = T625[3'h5:1'h0];
  assign T625 = T959 + 7'h1;
  assign T959 = {1'h0, R622};
  assign T626 = io_uarch_counters_12 != 1'h0;
  assign T960 = reset ? 58'h0 : T628;
  assign T628 = T630 ? T629 : R627;
  assign T629 = R627 + 58'h1;
  assign T630 = T626 & T631;
  assign T631 = T625[3'h6];
  assign T632 = T645 | T633;
  assign T633 = T133 ? T634 : 64'h0;
  assign T634 = {R640, R635};
  assign T961 = reset ? 6'h0 : T636;
  assign T636 = T639 ? T637 : R635;
  assign T637 = T638[3'h5:1'h0];
  assign T638 = T962 + 7'h1;
  assign T962 = {1'h0, R635};
  assign T639 = io_uarch_counters_11 != 1'h0;
  assign T963 = reset ? 58'h0 : T641;
  assign T641 = T643 ? T642 : R640;
  assign T642 = R640 + 58'h1;
  assign T643 = T639 & T644;
  assign T644 = T638[3'h6];
  assign T645 = T658 | T646;
  assign T646 = T135 ? T647 : 64'h0;
  assign T647 = {R653, R648};
  assign T964 = reset ? 6'h0 : T649;
  assign T649 = T652 ? T650 : R648;
  assign T650 = T651[3'h5:1'h0];
  assign T651 = T965 + 7'h1;
  assign T965 = {1'h0, R648};
  assign T652 = io_uarch_counters_10 != 1'h0;
  assign T966 = reset ? 58'h0 : T654;
  assign T654 = T656 ? T655 : R653;
  assign T655 = R653 + 58'h1;
  assign T656 = T652 & T657;
  assign T657 = T651[3'h6];
  assign T658 = T671 | T659;
  assign T659 = T137 ? T660 : 64'h0;
  assign T660 = {R666, R661};
  assign T967 = reset ? 6'h0 : T662;
  assign T662 = T665 ? T663 : R661;
  assign T663 = T664[3'h5:1'h0];
  assign T664 = T968 + 7'h1;
  assign T968 = {1'h0, R661};
  assign T665 = io_uarch_counters_9 != 1'h0;
  assign T969 = reset ? 58'h0 : T667;
  assign T667 = T669 ? T668 : R666;
  assign T668 = R666 + 58'h1;
  assign T669 = T665 & T670;
  assign T670 = T664[3'h6];
  assign T671 = T684 | T672;
  assign T672 = T139 ? T673 : 64'h0;
  assign T673 = {R679, R674};
  assign T970 = reset ? 6'h0 : T675;
  assign T675 = T678 ? T676 : R674;
  assign T676 = T677[3'h5:1'h0];
  assign T677 = T971 + 7'h1;
  assign T971 = {1'h0, R674};
  assign T678 = io_uarch_counters_8 != 1'h0;
  assign T972 = reset ? 58'h0 : T680;
  assign T680 = T682 ? T681 : R679;
  assign T681 = R679 + 58'h1;
  assign T682 = T678 & T683;
  assign T683 = T677[3'h6];
  assign T684 = T697 | T685;
  assign T685 = T141 ? T686 : 64'h0;
  assign T686 = {R692, R687};
  assign T973 = reset ? 6'h0 : T688;
  assign T688 = T691 ? T689 : R687;
  assign T689 = T690[3'h5:1'h0];
  assign T690 = T974 + 7'h1;
  assign T974 = {1'h0, R687};
  assign T691 = io_uarch_counters_7 != 1'h0;
  assign T975 = reset ? 58'h0 : T693;
  assign T693 = T695 ? T694 : R692;
  assign T694 = R692 + 58'h1;
  assign T695 = T691 & T696;
  assign T696 = T690[3'h6];
  assign T697 = T710 | T698;
  assign T698 = T143 ? T699 : 64'h0;
  assign T699 = {R705, R700};
  assign T976 = reset ? 6'h0 : T701;
  assign T701 = T704 ? T702 : R700;
  assign T702 = T703[3'h5:1'h0];
  assign T703 = T977 + 7'h1;
  assign T977 = {1'h0, R700};
  assign T704 = io_uarch_counters_6 != 1'h0;
  assign T978 = reset ? 58'h0 : T706;
  assign T706 = T708 ? T707 : R705;
  assign T707 = R705 + 58'h1;
  assign T708 = T704 & T709;
  assign T709 = T703[3'h6];
  assign T710 = T723 | T711;
  assign T711 = T145 ? T712 : 64'h0;
  assign T712 = {R718, R713};
  assign T979 = reset ? 6'h0 : T714;
  assign T714 = T717 ? T715 : R713;
  assign T715 = T716[3'h5:1'h0];
  assign T716 = T980 + 7'h1;
  assign T980 = {1'h0, R713};
  assign T717 = io_uarch_counters_5 != 1'h0;
  assign T981 = reset ? 58'h0 : T719;
  assign T719 = T721 ? T720 : R718;
  assign T720 = R718 + 58'h1;
  assign T721 = T717 & T722;
  assign T722 = T716[3'h6];
  assign T723 = T736 | T724;
  assign T724 = T147 ? T725 : 64'h0;
  assign T725 = {R731, R726};
  assign T982 = reset ? 6'h0 : T727;
  assign T727 = T730 ? T728 : R726;
  assign T728 = T729[3'h5:1'h0];
  assign T729 = T983 + 7'h1;
  assign T983 = {1'h0, R726};
  assign T730 = io_uarch_counters_4 != 1'h0;
  assign T984 = reset ? 58'h0 : T732;
  assign T732 = T734 ? T733 : R731;
  assign T733 = R731 + 58'h1;
  assign T734 = T730 & T735;
  assign T735 = T729[3'h6];
  assign T736 = T749 | T737;
  assign T737 = T149 ? T738 : 64'h0;
  assign T738 = {R744, R739};
  assign T985 = reset ? 6'h0 : T740;
  assign T740 = T743 ? T741 : R739;
  assign T741 = T742[3'h5:1'h0];
  assign T742 = T986 + 7'h1;
  assign T986 = {1'h0, R739};
  assign T743 = io_uarch_counters_3 != 1'h0;
  assign T987 = reset ? 58'h0 : T745;
  assign T745 = T747 ? T746 : R744;
  assign T746 = R744 + 58'h1;
  assign T747 = T743 & T748;
  assign T748 = T742[3'h6];
  assign T749 = T762 | T750;
  assign T750 = T151 ? T751 : 64'h0;
  assign T751 = {R757, R752};
  assign T988 = reset ? 6'h0 : T753;
  assign T753 = T756 ? T754 : R752;
  assign T754 = T755[3'h5:1'h0];
  assign T755 = T989 + 7'h1;
  assign T989 = {1'h0, R752};
  assign T756 = io_uarch_counters_2 != 1'h0;
  assign T990 = reset ? 58'h0 : T758;
  assign T758 = T760 ? T759 : R757;
  assign T759 = R757 + 58'h1;
  assign T760 = T756 & T761;
  assign T761 = T755[3'h6];
  assign T762 = T775 | T763;
  assign T763 = T153 ? T764 : 64'h0;
  assign T764 = {R770, R765};
  assign T991 = reset ? 6'h0 : T766;
  assign T766 = T769 ? T767 : R765;
  assign T767 = T768[3'h5:1'h0];
  assign T768 = T992 + 7'h1;
  assign T992 = {1'h0, R765};
  assign T769 = io_uarch_counters_1 != 1'h0;
  assign T993 = reset ? 58'h0 : T771;
  assign T771 = T773 ? T772 : R770;
  assign T772 = R770 + 58'h1;
  assign T773 = T769 & T774;
  assign T774 = T768[3'h6];
  assign T775 = T788 | T776;
  assign T776 = T155 ? T777 : 64'h0;
  assign T777 = {R783, R778};
  assign T994 = reset ? 6'h0 : T779;
  assign T779 = T782 ? T780 : R778;
  assign T780 = T781[3'h5:1'h0];
  assign T781 = T995 + 7'h1;
  assign T995 = {1'h0, R778};
  assign T782 = io_uarch_counters_0 != 1'h0;
  assign T996 = reset ? 58'h0 : T784;
  assign T784 = T786 ? T785 : R783;
  assign T785 = R783 + 58'h1;
  assign T786 = T782 & T787;
  assign T787 = T781[3'h6];
  assign T788 = T806 | T789;
  assign T789 = T157 ? T790 : 64'h0;
  assign T790 = {R799, R791};
  assign T997 = reset ? 6'h0 : T792;
  assign T792 = T798 ? T797 : T793;
  assign T793 = T796 ? T794 : R791;
  assign T794 = T795[3'h5:1'h0];
  assign T795 = T998 + 7'h1;
  assign T998 = {1'h0, R791};
  assign T796 = io_retire != 1'h0;
  assign T797 = wdata[3'h5:1'h0];
  assign T798 = wen & T157;
  assign T999 = reset ? 58'h0 : T800;
  assign T800 = T798 ? T805 : T801;
  assign T801 = T803 ? T802 : R799;
  assign T802 = R799 + 58'h1;
  assign T803 = T796 & T804;
  assign T804 = T795[3'h6];
  assign T805 = wdata[6'h3f:3'h6];
  assign T806 = T808 | T807;
  assign T807 = T159 ? T790 : 64'h0;
  assign T808 = T810 | T809;
  assign T809 = T161 ? reg_fromhost : 64'h0;
  assign T810 = T821 | T811;
  assign T811 = T163 ? reg_tohost : 64'h0;
  assign T1000 = reset ? 64'h0 : T812;
  assign T812 = T817 ? wdata : T813;
  assign T813 = T814 ? 64'h0 : reg_tohost;
  assign T814 = T815 & T163;
  assign T815 = host_csr_req_fire & T816;
  assign T816 = host_csr_bits_rw ^ 1'h1;
  assign T817 = T820 & T818;
  assign T818 = T819 | host_csr_req_fire;
  assign T819 = reg_tohost == 64'h0;
  assign T820 = wen & T163;
  assign T821 = T826 | T1001;
  assign T1001 = {63'h0, T822};
  assign T822 = T165 ? reg_stats : 1'h0;
  assign T1002 = reset ? 1'h0 : T823;
  assign T823 = T825 ? T824 : reg_stats;
  assign T824 = wdata[1'h0];
  assign T825 = wen & T165;
  assign T826 = T828 | T1003;
  assign T1003 = {63'h0, T827};
  assign T827 = T167 ? io_host_id : 1'h0;
  assign T828 = T830 | T829;
  assign T829 = T169 ? reg_mtimecmp : 64'h0;
  assign T830 = T832 | T831;
  assign T831 = T171 ? reg_mcause : 64'h0;
  assign T832 = T837 | T833;
  assign T833 = T173 ? T834 : 64'h0;
  assign T834 = {T835, reg_mbadaddr};
  assign T835 = 24'h0 - T1004;
  assign T1004 = {23'h0, T836};
  assign T836 = reg_mbadaddr[6'h27];
  assign T837 = T842 | T838;
  assign T838 = T175 ? T839 : 64'h0;
  assign T839 = {T840, reg_mepc};
  assign T840 = 24'h0 - T1005;
  assign T1005 = {23'h0, T841};
  assign T841 = reg_mepc[6'h27];
  assign T842 = T846 | T843;
  assign T843 = T177 ? reg_mscratch : 64'h0;
  assign T844 = T845 ? wdata : reg_mscratch;
  assign T845 = wen & T177;
  assign T846 = T856 | T1006;
  assign T1006 = {56'h0, T847};
  assign T847 = T179 ? T848 : 8'h0;
  assign T848 = T849;
  assign T849 = {T853, T850};
  assign T850 = {T852, T851};
  assign T851 = {reg_mie_ssip, reg_mie_usip};
  assign T1007 = reset ? 1'h0 : reg_mie_usip;
  assign T852 = {reg_mie_msip, reg_mie_hsip};
  assign T1008 = reset ? 1'h0 : reg_mie_hsip;
  assign T853 = {T855, T854};
  assign T854 = {reg_mie_stip, reg_mie_utip};
  assign T1009 = reset ? 1'h0 : reg_mie_utip;
  assign T855 = {reg_mie_mtip, reg_mie_htip};
  assign T1010 = reset ? 1'h0 : reg_mie_htip;
  assign T856 = T866 | T1011;
  assign T1011 = {56'h0, T857};
  assign T857 = T181 ? T858 : 8'h0;
  assign T858 = T859;
  assign T859 = {T863, T860};
  assign T860 = {T862, T861};
  assign T861 = {reg_mip_ssip, reg_mip_usip};
  assign T1012 = reset ? 1'h0 : reg_mip_usip;
  assign T862 = {reg_mip_msip, reg_mip_hsip};
  assign T1013 = reset ? 1'h0 : reg_mip_hsip;
  assign T863 = {T865, T864};
  assign T864 = {reg_mip_stip, reg_mip_utip};
  assign T1014 = reset ? 1'h0 : reg_mip_utip;
  assign T865 = {reg_mip_mtip, reg_mip_htip};
  assign T1015 = reset ? 1'h0 : reg_mip_htip;
  assign T866 = T867 | 64'h0;
  assign T867 = T869 | T1016;
  assign T1016 = {33'h0, T868};
  assign T868 = T185 ? 31'h40000000 : 31'h0;
  assign T869 = T871 | T870;
  assign T870 = T187 ? reg_mtvec : 64'h0;
  assign T871 = T872 | 64'h0;
  assign T872 = T873 | 64'h0;
  assign T873 = T875 | T874;
  assign T874 = T59 ? read_mstatus : 64'h0;
  assign T875 = T876 | T1017;
  assign T1017 = {63'h0, T194};
  assign T876 = T878 | T877;
  assign T877 = T196 ? 64'h8000000000841129 : 64'h0;
  assign T878 = T880 | T879;
  assign T879 = T198 ? read_time : 64'h0;
  assign T880 = T882 | T881;
  assign T881 = T200 ? read_time : 64'h0;
  assign T882 = T884 | T883;
  assign T883 = T202 ? read_time : 64'h0;
  assign T884 = T886 | T885;
  assign T885 = T204 ? read_time : 64'h0;
  assign T886 = T888 | T887;
  assign T887 = T206 ? read_time : 64'h0;
  assign T888 = T890 | T889;
  assign T889 = T208 ? T323 : 64'h0;
  assign T890 = T1018 | T891;
  assign T891 = T210 ? T323 : 64'h0;
  assign T1018 = {56'h0, T892};
  assign T892 = T1021 | T893;
  assign T893 = T100 ? T894 : 8'h0;
  assign T894 = {reg_frm, reg_fflags};
  assign T1019 = T895[3'h4:1'h0];
  assign T895 = T322 ? wdata : T896;
  assign T896 = T899 ? wdata : T1020;
  assign T1020 = {59'h0, T897};
  assign T897 = io_fcsr_flags_valid ? T898 : reg_fflags;
  assign T898 = reg_fflags | io_fcsr_flags_bits;
  assign T899 = wen & T103;
  assign T1021 = {3'h0, T900};
  assign T900 = T902 | T1022;
  assign T1022 = {2'h0, T901};
  assign T901 = T102 ? reg_frm : 3'h0;
  assign T902 = T103 ? reg_fflags : 5'h0;
  assign io_host_debug_stats_csr = reg_stats;
  assign io_host_csr_resp_bits = host_csr_bits_data;
  assign io_host_csr_resp_valid = host_csr_rep_valid;
  assign T903 = T905 ? 1'h0 : T904;
  assign T904 = host_csr_req_fire ? 1'h1 : host_csr_rep_valid;
  assign T905 = io_host_csr_resp_ready & io_host_csr_resp_valid;
  assign io_host_csr_req_ready = T906;
  assign T906 = T908 & T907;
  assign T907 = host_csr_rep_valid ^ 1'h1;
  assign T908 = host_csr_req_valid ^ 1'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "these conditions must be mutually exclusive");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if(T88) begin
      reg_mstatus_prv <= T87;
    end else if(insn_redirect_trap) begin
      reg_mstatus_prv <= 2'h1;
    end else if(insn_ret) begin
      reg_mstatus_prv <= reg_mstatus_prv1;
    end else if(T25) begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_prv1 <= 2'h3;
    end else if(T76) begin
      reg_mstatus_prv1 <= T909;
    end else if(T69) begin
      reg_mstatus_prv1 <= T68;
    end else if(insn_ret) begin
      reg_mstatus_prv1 <= reg_mstatus_prv2;
    end else if(T25) begin
      reg_mstatus_prv1 <= reg_mstatus_prv;
    end
    if(reset) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T52) begin
      reg_mstatus_prv2 <= T35;
    end else if(insn_ret) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T25) begin
      reg_mstatus_prv2 <= reg_mstatus_prv1;
    end
    if(host_csr_req_fire) begin
      host_csr_bits_data <= io_rw_rdata;
    end else if(T40) begin
      host_csr_bits_data <= io_host_csr_req_bits_data;
    end
    if(host_csr_req_fire) begin
      host_csr_req_valid <= 1'h0;
    end else if(T40) begin
      host_csr_req_valid <= 1'h1;
    end
    if(T40) begin
      host_csr_bits_addr <= io_host_csr_req_bits_addr;
    end
    if(T40) begin
      host_csr_bits_rw <= io_host_csr_req_bits_rw;
    end
    if(reset) begin
      reg_mstatus_ie <= 1'h0;
    end else if(T76) begin
      reg_mstatus_ie <= T244;
    end else if(T58) begin
      reg_mstatus_ie <= T243;
    end else if(insn_ret) begin
      reg_mstatus_ie <= reg_mstatus_ie1;
    end else if(T25) begin
      reg_mstatus_ie <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_ie1 <= 1'h0;
    end else if(T76) begin
      reg_mstatus_ie1 <= T242;
    end else if(T58) begin
      reg_mstatus_ie1 <= T241;
    end else if(insn_ret) begin
      reg_mstatus_ie1 <= reg_mstatus_ie2;
    end else if(T25) begin
      reg_mstatus_ie1 <= reg_mstatus_ie;
    end
    if(reset) begin
      reg_mstatus_ie2 <= 1'h0;
    end else if(T58) begin
      reg_mstatus_ie2 <= T240;
    end else if(insn_ret) begin
      reg_mstatus_ie2 <= 1'h1;
    end else if(T25) begin
      reg_mstatus_ie2 <= reg_mstatus_ie1;
    end
    if(reset) begin
      reg_mip_ssip <= 1'h0;
    end else if(T253) begin
      reg_mip_ssip <= T252;
    end else if(T251) begin
      reg_mip_ssip <= T250;
    end
    if(reset) begin
      reg_mie_ssip <= 1'h0;
    end else if(T259) begin
      reg_mie_ssip <= T258;
    end else if(T257) begin
      reg_mie_ssip <= T256;
    end
    if(reset) begin
      reg_mip_msip <= 1'h0;
    end else if(T270) begin
      reg_mip_msip <= T269;
    end else if(T251) begin
      reg_mip_msip <= T268;
    end
    if(reset) begin
      reg_mie_msip <= 1'h0;
    end else if(T257) begin
      reg_mie_msip <= T272;
    end
    if(reset) begin
      reg_mip_stip <= 1'h0;
    end else if(T251) begin
      reg_mip_stip <= T280;
    end
    if(reset) begin
      reg_mie_stip <= 1'h0;
    end else if(T259) begin
      reg_mie_stip <= T284;
    end else if(T257) begin
      reg_mie_stip <= T283;
    end
    if(reset) begin
      reg_mip_mtip <= 1'h0;
    end else if(T297) begin
      reg_mip_mtip <= 1'h0;
    end else if(T293) begin
      reg_mip_mtip <= 1'h1;
    end
    if(T295) begin
      read_time <= wdata;
    end
    if(T297) begin
      reg_mtimecmp <= wdata;
    end
    if(reset) begin
      reg_mie_mtip <= 1'h0;
    end else if(T257) begin
      reg_mie_mtip <= T299;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T307) begin
      reg_fromhost <= wdata;
    end
    reg_frm <= T922;
    if(reset) begin
      R324 <= 6'h0;
    end else begin
      R324 <= T325;
    end
    if(reset) begin
      R327 <= 58'h0;
    end else if(T330) begin
      R327 <= T329;
    end
    reg_sepc <= T930;
    reg_mepc <= T932;
    reg_stvec <= T934;
    if(reset) begin
      reg_mtvec <= 64'h100;
    end else if(T367) begin
      reg_mtvec <= T366;
    end
    if(T373) begin
      reg_sptbr <= T371;
    end
    if(reset) begin
      reg_mstatus_ie3 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_prv3 <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if(T76) begin
      reg_mstatus_fs <= T382;
    end else if(T58) begin
      reg_mstatus_fs <= T381;
    end
    if(reset) begin
      reg_mstatus_xs <= 2'h0;
    end else if(T76) begin
      reg_mstatus_xs <= T389;
    end else if(T58) begin
      reg_mstatus_xs <= T388;
    end
    if(reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if(T76) begin
      reg_mstatus_mprv <= T395;
    end else if(T58) begin
      reg_mstatus_mprv <= T394;
    end else if(T25) begin
      reg_mstatus_mprv <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_vm <= 5'h0;
    end else if(T402) begin
      reg_mstatus_vm <= 5'h9;
    end else if(T399) begin
      reg_mstatus_vm <= 5'h0;
    end
    if(reset) begin
      reg_mstatus_zero1 <= 9'h0;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_zero2 <= 31'h0;
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else if(some_interrupt_pending) begin
      reg_wfi <= 1'h0;
    end else if(insn_wfi) begin
      reg_wfi <= 1'h1;
    end
    if(insn_redirect_trap) begin
      reg_sbadaddr <= reg_mbadaddr;
    end
    if(T474) begin
      reg_mbadaddr <= T473;
    end else if(T465) begin
      reg_mbadaddr <= T457;
    end else if(T25) begin
      reg_mbadaddr <= io_pc;
    end
    if(insn_redirect_trap) begin
      reg_scause <= reg_mcause;
    end
    if(T490) begin
      reg_mcause <= T489;
    end else if(T488) begin
      reg_mcause <= T945;
    end else if(T486) begin
      reg_mcause <= 64'h3;
    end else if(T485) begin
      reg_mcause <= 64'h2;
    end else if(T25) begin
      reg_mcause <= io_cause;
    end
    if(T494) begin
      reg_sscratch <= wdata;
    end
    if(reset) begin
      R583 <= 6'h0;
    end else if(T587) begin
      R583 <= T585;
    end
    if(reset) begin
      R588 <= 58'h0;
    end else if(T591) begin
      R588 <= T590;
    end
    if(reset) begin
      R596 <= 6'h0;
    end else if(T600) begin
      R596 <= T598;
    end
    if(reset) begin
      R601 <= 58'h0;
    end else if(T604) begin
      R601 <= T603;
    end
    if(reset) begin
      R609 <= 6'h0;
    end else if(T613) begin
      R609 <= T611;
    end
    if(reset) begin
      R614 <= 58'h0;
    end else if(T617) begin
      R614 <= T616;
    end
    if(reset) begin
      R622 <= 6'h0;
    end else if(T626) begin
      R622 <= T624;
    end
    if(reset) begin
      R627 <= 58'h0;
    end else if(T630) begin
      R627 <= T629;
    end
    if(reset) begin
      R635 <= 6'h0;
    end else if(T639) begin
      R635 <= T637;
    end
    if(reset) begin
      R640 <= 58'h0;
    end else if(T643) begin
      R640 <= T642;
    end
    if(reset) begin
      R648 <= 6'h0;
    end else if(T652) begin
      R648 <= T650;
    end
    if(reset) begin
      R653 <= 58'h0;
    end else if(T656) begin
      R653 <= T655;
    end
    if(reset) begin
      R661 <= 6'h0;
    end else if(T665) begin
      R661 <= T663;
    end
    if(reset) begin
      R666 <= 58'h0;
    end else if(T669) begin
      R666 <= T668;
    end
    if(reset) begin
      R674 <= 6'h0;
    end else if(T678) begin
      R674 <= T676;
    end
    if(reset) begin
      R679 <= 58'h0;
    end else if(T682) begin
      R679 <= T681;
    end
    if(reset) begin
      R687 <= 6'h0;
    end else if(T691) begin
      R687 <= T689;
    end
    if(reset) begin
      R692 <= 58'h0;
    end else if(T695) begin
      R692 <= T694;
    end
    if(reset) begin
      R700 <= 6'h0;
    end else if(T704) begin
      R700 <= T702;
    end
    if(reset) begin
      R705 <= 58'h0;
    end else if(T708) begin
      R705 <= T707;
    end
    if(reset) begin
      R713 <= 6'h0;
    end else if(T717) begin
      R713 <= T715;
    end
    if(reset) begin
      R718 <= 58'h0;
    end else if(T721) begin
      R718 <= T720;
    end
    if(reset) begin
      R726 <= 6'h0;
    end else if(T730) begin
      R726 <= T728;
    end
    if(reset) begin
      R731 <= 58'h0;
    end else if(T734) begin
      R731 <= T733;
    end
    if(reset) begin
      R739 <= 6'h0;
    end else if(T743) begin
      R739 <= T741;
    end
    if(reset) begin
      R744 <= 58'h0;
    end else if(T747) begin
      R744 <= T746;
    end
    if(reset) begin
      R752 <= 6'h0;
    end else if(T756) begin
      R752 <= T754;
    end
    if(reset) begin
      R757 <= 58'h0;
    end else if(T760) begin
      R757 <= T759;
    end
    if(reset) begin
      R765 <= 6'h0;
    end else if(T769) begin
      R765 <= T767;
    end
    if(reset) begin
      R770 <= 58'h0;
    end else if(T773) begin
      R770 <= T772;
    end
    if(reset) begin
      R778 <= 6'h0;
    end else if(T782) begin
      R778 <= T780;
    end
    if(reset) begin
      R783 <= 58'h0;
    end else if(T786) begin
      R783 <= T785;
    end
    if(reset) begin
      R791 <= 6'h0;
    end else if(T798) begin
      R791 <= T797;
    end else if(T796) begin
      R791 <= T794;
    end
    if(reset) begin
      R799 <= 58'h0;
    end else if(T798) begin
      R799 <= T805;
    end else if(T803) begin
      R799 <= T802;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T817) begin
      reg_tohost <= wdata;
    end else if(T814) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T825) begin
      reg_stats <= T824;
    end
    if(T845) begin
      reg_mscratch <= wdata;
    end
    if(reset) begin
      reg_mie_usip <= 1'h0;
    end
    if(reset) begin
      reg_mie_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mie_utip <= 1'h0;
    end
    if(reset) begin
      reg_mie_htip <= 1'h0;
    end
    if(reset) begin
      reg_mip_usip <= 1'h0;
    end
    if(reset) begin
      reg_mip_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mip_utip <= 1'h0;
    end
    if(reset) begin
      reg_mip_htip <= 1'h0;
    end
    reg_fflags <= T1019;
    if(T905) begin
      host_csr_rep_valid <= 1'h0;
    end else if(host_csr_req_fire) begin
      host_csr_rep_valid <= 1'h1;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out,
    output io_cmp_out
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[63:0] in1_xor_in2;
  wire[63:0] in2_inv;
  wire[63:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[63:0] T17;
  wire[63:0] T146;
  wire T18;
  wire[63:0] T19;
  wire[63:0] T20;
  wire[63:0] out;
  wire[63:0] shift_logic;
  wire[63:0] shout;
  wire[63:0] T21;
  wire[63:0] shout_l;
  wire[63:0] T22;
  wire[63:0] T23;
  wire[62:0] T24;
  wire[63:0] T25;
  wire[63:0] T26;
  wire[63:0] T27;
  wire[61:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] T31;
  wire[59:0] T32;
  wire[63:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[55:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[47:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[31:0] T44;
  wire[63:0] shout_r;
  wire[64:0] T45;
  wire[5:0] shamt;
  wire[4:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[64:0] T51;
  wire[64:0] T52;
  wire[63:0] shin;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] T55;
  wire[62:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[61:0] T60;
  wire[63:0] T61;
  wire[63:0] T62;
  wire[63:0] T63;
  wire[59:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire[63:0] T67;
  wire[55:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire[47:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  wire[31:0] T76;
  wire[63:0] T77;
  wire[63:0] T147;
  wire[31:0] T78;
  wire[63:0] T79;
  wire[63:0] T148;
  wire[47:0] T80;
  wire[63:0] T81;
  wire[63:0] T149;
  wire[55:0] T82;
  wire[63:0] T83;
  wire[63:0] T150;
  wire[59:0] T84;
  wire[63:0] T85;
  wire[63:0] T151;
  wire[61:0] T86;
  wire[63:0] T87;
  wire[63:0] T152;
  wire[62:0] T88;
  wire[63:0] shin_r;
  wire[31:0] T89;
  wire[31:0] T90;
  wire[31:0] T91;
  wire[31:0] T153;
  wire T92;
  wire T93;
  wire T94;
  wire[31:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[63:0] T104;
  wire[63:0] T154;
  wire[31:0] T105;
  wire[63:0] T106;
  wire[63:0] T155;
  wire[47:0] T107;
  wire[63:0] T108;
  wire[63:0] T156;
  wire[55:0] T109;
  wire[63:0] T110;
  wire[63:0] T157;
  wire[59:0] T111;
  wire[63:0] T112;
  wire[63:0] T158;
  wire[61:0] T113;
  wire[63:0] T114;
  wire[63:0] T159;
  wire[62:0] T115;
  wire T116;
  wire[63:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire[63:0] T121;
  wire[63:0] logic;
  wire[63:0] T122;
  wire[63:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[63:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[63:0] T160;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[63:0] T140;
  wire[31:0] T141;
  wire[31:0] T142;
  wire[31:0] T161;
  wire T143;
  wire T144;
  wire T145;


  assign io_cmp_out = T0;
  assign T0 = T16 ^ T1;
  assign T1 = T14 ? T11 : T2;
  assign T2 = T8 ? T7 : T3;
  assign T3 = T6 ? T5 : T4;
  assign T4 = io_in1[6'h3f];
  assign T5 = io_in2[6'h3f];
  assign T6 = io_fn[1'h1];
  assign T7 = io_adder_out[6'h3f];
  assign T8 = T10 == T9;
  assign T9 = io_in2[6'h3f];
  assign T10 = io_in1[6'h3f];
  assign T11 = in1_xor_in2 == 64'h0;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign in2_inv = T13 ? T12 : io_in2;
  assign T12 = ~ io_in2;
  assign T13 = io_fn[2'h3];
  assign T14 = T15 ^ 1'h1;
  assign T15 = io_fn[2'h3];
  assign T16 = io_fn[1'h0];
  assign io_adder_out = T17;
  assign T17 = T19 + T146;
  assign T146 = {63'h0, T18};
  assign T18 = io_fn[2'h3];
  assign T19 = io_in1 + in2_inv;
  assign io_out = T20;
  assign T20 = T144 ? T140 : out;
  assign out = T137 ? io_adder_out : shift_logic;
  assign shift_logic = T121 | shout;
  assign shout = T117 | T21;
  assign T21 = T116 ? shout_l : 64'h0;
  assign shout_l = T114 | T22;
  assign T22 = T23 & 64'haaaaaaaaaaaaaaaa;
  assign T23 = T24 << 1'h1;
  assign T24 = T25[6'h3e:1'h0];
  assign T25 = T112 | T26;
  assign T26 = T27 & 64'hcccccccccccccccc;
  assign T27 = T28 << 2'h2;
  assign T28 = T29[6'h3d:1'h0];
  assign T29 = T110 | T30;
  assign T30 = T31 & 64'hf0f0f0f0f0f0f0f0;
  assign T31 = T32 << 3'h4;
  assign T32 = T33[6'h3b:1'h0];
  assign T33 = T108 | T34;
  assign T34 = T35 & 64'hff00ff00ff00ff00;
  assign T35 = T36 << 4'h8;
  assign T36 = T37[6'h37:1'h0];
  assign T37 = T106 | T38;
  assign T38 = T39 & 64'hffff0000ffff0000;
  assign T39 = T40 << 5'h10;
  assign T40 = T41[6'h2f:1'h0];
  assign T41 = T104 | T42;
  assign T42 = T43 & 64'hffffffff00000000;
  assign T43 = T44 << 6'h20;
  assign T44 = shout_r[5'h1f:1'h0];
  assign shout_r = T45[6'h3f:1'h0];
  assign T45 = $signed(T51) >>> shamt;
  assign shamt = {T47, T46};
  assign T46 = io_in2[3'h4:1'h0];
  assign T47 = T50 & T48;
  assign T48 = 1'h1 == T49;
  assign T49 = io_dw & 1'h1;
  assign T50 = io_in2[3'h5];
  assign T51 = T52;
  assign T52 = {T101, shin};
  assign shin = T98 ? shin_r : T53;
  assign T53 = T87 | T54;
  assign T54 = T55 & 64'haaaaaaaaaaaaaaaa;
  assign T55 = T56 << 1'h1;
  assign T56 = T57[6'h3e:1'h0];
  assign T57 = T85 | T58;
  assign T58 = T59 & 64'hcccccccccccccccc;
  assign T59 = T60 << 2'h2;
  assign T60 = T61[6'h3d:1'h0];
  assign T61 = T83 | T62;
  assign T62 = T63 & 64'hf0f0f0f0f0f0f0f0;
  assign T63 = T64 << 3'h4;
  assign T64 = T65[6'h3b:1'h0];
  assign T65 = T81 | T66;
  assign T66 = T67 & 64'hff00ff00ff00ff00;
  assign T67 = T68 << 4'h8;
  assign T68 = T69[6'h37:1'h0];
  assign T69 = T79 | T70;
  assign T70 = T71 & 64'hffff0000ffff0000;
  assign T71 = T72 << 5'h10;
  assign T72 = T73[6'h2f:1'h0];
  assign T73 = T77 | T74;
  assign T74 = T75 & 64'hffffffff00000000;
  assign T75 = T76 << 6'h20;
  assign T76 = shin_r[5'h1f:1'h0];
  assign T77 = T147 & 64'hffffffff;
  assign T147 = {32'h0, T78};
  assign T78 = shin_r >> 6'h20;
  assign T79 = T148 & 64'hffff0000ffff;
  assign T148 = {16'h0, T80};
  assign T80 = T73 >> 5'h10;
  assign T81 = T149 & 64'hff00ff00ff00ff;
  assign T149 = {8'h0, T82};
  assign T82 = T69 >> 4'h8;
  assign T83 = T150 & 64'hf0f0f0f0f0f0f0f;
  assign T150 = {4'h0, T84};
  assign T84 = T65 >> 3'h4;
  assign T85 = T151 & 64'h3333333333333333;
  assign T151 = {2'h0, T86};
  assign T86 = T61 >> 2'h2;
  assign T87 = T152 & 64'h5555555555555555;
  assign T152 = {1'h0, T88};
  assign T88 = T57 >> 1'h1;
  assign shin_r = {T90, T89};
  assign T89 = io_in1[5'h1f:1'h0];
  assign T90 = T96 ? T95 : T91;
  assign T91 = 32'h0 - T153;
  assign T153 = {31'h0, T92};
  assign T92 = T94 & T93;
  assign T93 = io_in1[5'h1f];
  assign T94 = io_fn[2'h3];
  assign T95 = io_in1[6'h3f:6'h20];
  assign T96 = 1'h1 == T97;
  assign T97 = io_dw & 1'h1;
  assign T98 = T100 | T99;
  assign T99 = io_fn == 4'hb;
  assign T100 = io_fn == 4'h5;
  assign T101 = T103 & T102;
  assign T102 = shin[6'h3f];
  assign T103 = io_fn[2'h3];
  assign T104 = T154 & 64'hffffffff;
  assign T154 = {32'h0, T105};
  assign T105 = shout_r >> 6'h20;
  assign T106 = T155 & 64'hffff0000ffff;
  assign T155 = {16'h0, T107};
  assign T107 = T41 >> 5'h10;
  assign T108 = T156 & 64'hff00ff00ff00ff;
  assign T156 = {8'h0, T109};
  assign T109 = T37 >> 4'h8;
  assign T110 = T157 & 64'hf0f0f0f0f0f0f0f;
  assign T157 = {4'h0, T111};
  assign T111 = T33 >> 3'h4;
  assign T112 = T158 & 64'h3333333333333333;
  assign T158 = {2'h0, T113};
  assign T113 = T29 >> 2'h2;
  assign T114 = T159 & 64'h5555555555555555;
  assign T159 = {1'h0, T115};
  assign T115 = T25 >> 1'h1;
  assign T116 = io_fn == 4'h1;
  assign T117 = T118 ? shout_r : 64'h0;
  assign T118 = T120 | T119;
  assign T119 = io_fn == 4'hb;
  assign T120 = io_fn == 4'h5;
  assign T121 = T160 | logic;
  assign logic = T127 | T122;
  assign T122 = T124 ? T123 : 64'h0;
  assign T123 = io_in1 & io_in2;
  assign T124 = T126 | T125;
  assign T125 = io_fn == 4'h7;
  assign T126 = io_fn == 4'h6;
  assign T127 = T128 ? in1_xor_in2 : 64'h0;
  assign T128 = T130 | T129;
  assign T129 = io_fn == 4'h6;
  assign T130 = io_fn == 4'h4;
  assign T160 = {63'h0, T131};
  assign T131 = T132 & io_cmp_out;
  assign T132 = T134 | T133;
  assign T133 = 4'hc <= io_fn;
  assign T134 = T136 | T135;
  assign T135 = io_fn == 4'h3;
  assign T136 = io_fn == 4'h2;
  assign T137 = T139 | T138;
  assign T138 = io_fn == 4'ha;
  assign T139 = io_fn == 4'h0;
  assign T140 = {T142, T141};
  assign T141 = out[5'h1f:1'h0];
  assign T142 = 32'h0 - T161;
  assign T161 = {31'h0, T143};
  assign T143 = out[5'h1f];
  assign T144 = 1'h0 == T145;
  assign T145 = io_dw & 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[129:0] T188;
  wire[63:0] negated_remainder;
  wire[63:0] T126;
  wire T11;
  wire T12;
  reg  isMul;
  wire T13;
  wire cmdMul;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  reg [2:0] state;
  wire[2:0] T189;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  reg  neg_out;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  isHi;
  wire T34;
  wire cmdHi;
  wire T35;
  wire T36;
  wire T37;
  wire[3:0] T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T43;
  wire[64:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[64:0] T48;
  wire[63:0] rhs_in;
  wire[31:0] T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] T190;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire rhs_sign;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire rhsSigned;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire[64:0] T63;
  wire T64;
  reg [6:0] count;
  wire[6:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[6:0] T68;
  wire[6:0] T69;
  wire[6:0] T70;
  wire[6:0] T191;
  wire[5:0] T71;
  wire[5:0] T72;
  wire[5:0] T73;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[5:0] T221;
  wire[5:0] T222;
  wire[5:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire[4:0] T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire[4:0] T231;
  wire[4:0] T232;
  wire[4:0] T233;
  wire[4:0] T234;
  wire[4:0] T235;
  wire[4:0] T236;
  wire[4:0] T237;
  wire[4:0] T238;
  wire[4:0] T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[3:0] T246;
  wire[3:0] T247;
  wire[2:0] T248;
  wire[2:0] T249;
  wire[2:0] T250;
  wire[2:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire T254;
  wire[63:0] T75;
  wire[63:0] T76;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire[5:0] T77;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[5:0] T321;
  wire[5:0] T322;
  wire[5:0] T323;
  wire[5:0] T324;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[5:0] T329;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[4:0] T357;
  wire[4:0] T358;
  wire[4:0] T359;
  wire[4:0] T360;
  wire[4:0] T361;
  wire[4:0] T362;
  wire[4:0] T363;
  wire[4:0] T364;
  wire[3:0] T365;
  wire[3:0] T366;
  wire[3:0] T367;
  wire[3:0] T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[2:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire[2:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire T379;
  wire[63:0] T79;
  wire[63:0] T80;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire lhs_sign;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire lhsSigned;
  wire T90;
  wire T91;
  wire[3:0] T92;
  wire T93;
  wire T94;
  wire[2:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[63:0] T103;
  wire[64:0] T104;
  wire[5:0] T105;
  wire[10:0] T106;
  wire[63:0] T107;
  wire[128:0] T108;
  wire[63:0] T109;
  wire[64:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire[129:0] T442;
  wire T127;
  wire[129:0] T443;
  wire[63:0] T128;
  wire T129;
  wire[129:0] T130;
  wire[64:0] T131;
  wire[63:0] T132;
  wire[128:0] T133;
  wire[63:0] T134;
  wire[128:0] T135;
  wire[128:0] T136;
  wire[128:0] T137;
  wire[55:0] T138;
  wire[72:0] T139;
  wire[72:0] T444;
  wire[64:0] T140;
  wire[64:0] T141;
  wire[7:0] T445;
  wire T446;
  wire[72:0] T142;
  wire[8:0] T143;
  wire[8:0] T144;
  wire[7:0] T145;
  wire[64:0] T146;
  wire[128:0] T147;
  wire[5:0] T148;
  wire[10:0] T149;
  wire[10:0] T150;
  wire[64:0] T151;
  wire[64:0] T152;
  wire T153;
  wire T154;
  wire[129:0] T447;
  wire[128:0] T155;
  wire[64:0] T156;
  wire T157;
  wire[63:0] T158;
  wire[63:0] T159;
  wire[63:0] T160;
  wire[63:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire[129:0] T448;
  wire[126:0] T165;
  wire[63:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[129:0] T449;
  wire[63:0] lhs_in;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T450;
  wire[31:0] T176;
  wire T177;
  wire T178;
  wire[63:0] T179;
  wire[31:0] T180;
  wire[31:0] T181;
  wire[31:0] T451;
  wire T182;
  wire T183;
  wire T184;
  reg  req_dw;
  wire T185;
  wire T186;
  wire T187;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T183 ? T179 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T449 : T5;
  assign T5 = T167 ? T448 : T6;
  assign T6 = T162 ? T447 : T7;
  assign T7 = T153 ? T130 : T8;
  assign T8 = T129 ? T443 : T9;
  assign T9 = T127 ? T442 : T10;
  assign T10 = T11 ? T188 : remainder;
  assign T188 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T126;
  assign T126 = remainder[6'h3f:1'h0];
  assign T11 = T20 & T12;
  assign T12 = T19 | isMul;
  assign T13 = T1 ? cmdMul : isMul;
  assign cmdMul = T14;
  assign T14 = T17 | T15;
  assign T15 = T16 == 4'h8;
  assign T16 = io_req_bits_fn & 4'h8;
  assign T17 = T18 == 4'h0;
  assign T18 = io_req_bits_fn & 4'h4;
  assign T19 = remainder[6'h3f];
  assign T20 = state == 3'h1;
  assign T189 = reset ? 3'h0 : T21;
  assign T21 = T1 ? T122 : T22;
  assign T22 = T120 ? 3'h0 : T23;
  assign T23 = T118 ? T116 : T24;
  assign T24 = T96 ? T95 : T25;
  assign T25 = T129 ? T28 : T26;
  assign T26 = T127 ? 3'h5 : T27;
  assign T27 = T20 ? 3'h2 : state;
  assign T28 = neg_out ? 3'h4 : 3'h5;
  assign T29 = T1 ? T82 : T30;
  assign T30 = T31 ? 1'h0 : neg_out;
  assign T31 = T162 & T32;
  assign T32 = T41 & T33;
  assign T33 = isHi ^ 1'h1;
  assign T34 = T1 ? cmdHi : isHi;
  assign cmdHi = T35;
  assign T35 = T36 | T15;
  assign T36 = T39 | T37;
  assign T37 = T38 == 4'h2;
  assign T38 = io_req_bits_fn & 4'h2;
  assign T39 = T40 == 4'h1;
  assign T40 = io_req_bits_fn & 4'h5;
  assign T41 = T64 & T42;
  assign T42 = less ^ 1'h1;
  assign less = subtractor[7'h40];
  assign subtractor = T63 - divisor;
  assign T43 = T1 ? T48 : T44;
  assign T44 = T45 ? subtractor : divisor;
  assign T45 = T20 & T46;
  assign T46 = T47 | isMul;
  assign T47 = divisor[6'h3f];
  assign T48 = {rhs_sign, rhs_in};
  assign rhs_in = {T50, T49};
  assign T49 = io_req_bits_in2[5'h1f:1'h0];
  assign T50 = T53 ? T52 : T51;
  assign T51 = 32'h0 - T190;
  assign T190 = {31'h0, rhs_sign};
  assign T52 = io_req_bits_in2[6'h3f:6'h20];
  assign T53 = 1'h1 == T54;
  assign T54 = io_req_bits_dw & 1'h1;
  assign rhs_sign = rhsSigned & T55;
  assign T55 = T58 ? T57 : T56;
  assign T56 = io_req_bits_in2[5'h1f];
  assign T57 = io_req_bits_in2[6'h3f];
  assign T58 = 1'h1 == T59;
  assign T59 = io_req_bits_dw & 1'h1;
  assign rhsSigned = T60;
  assign T60 = T61 | T17;
  assign T61 = T62 == 4'h0;
  assign T62 = io_req_bits_fn & 4'h9;
  assign T63 = remainder[8'h80:7'h40];
  assign T64 = count == 7'h0;
  assign T65 = T1 ? 7'h0 : T66;
  assign T66 = T167 ? T191 : T67;
  assign T67 = T162 ? T70 : T68;
  assign T68 = T153 ? T69 : count;
  assign T69 = count + 7'h1;
  assign T70 = count + 7'h1;
  assign T191 = {1'h0, T71};
  assign T71 = T81 ? 6'h3f : T72;
  assign T72 = T73;
  assign T73 = T77 - T192;
  assign T192 = T316 ? 6'h3f : T193;
  assign T193 = T315 ? 6'h3e : T194;
  assign T194 = T314 ? 6'h3d : T195;
  assign T195 = T313 ? 6'h3c : T196;
  assign T196 = T312 ? 6'h3b : T197;
  assign T197 = T311 ? 6'h3a : T198;
  assign T198 = T310 ? 6'h39 : T199;
  assign T199 = T309 ? 6'h38 : T200;
  assign T200 = T308 ? 6'h37 : T201;
  assign T201 = T307 ? 6'h36 : T202;
  assign T202 = T306 ? 6'h35 : T203;
  assign T203 = T305 ? 6'h34 : T204;
  assign T204 = T304 ? 6'h33 : T205;
  assign T205 = T303 ? 6'h32 : T206;
  assign T206 = T302 ? 6'h31 : T207;
  assign T207 = T301 ? 6'h30 : T208;
  assign T208 = T300 ? 6'h2f : T209;
  assign T209 = T299 ? 6'h2e : T210;
  assign T210 = T298 ? 6'h2d : T211;
  assign T211 = T297 ? 6'h2c : T212;
  assign T212 = T296 ? 6'h2b : T213;
  assign T213 = T295 ? 6'h2a : T214;
  assign T214 = T294 ? 6'h29 : T215;
  assign T215 = T293 ? 6'h28 : T216;
  assign T216 = T292 ? 6'h27 : T217;
  assign T217 = T291 ? 6'h26 : T218;
  assign T218 = T290 ? 6'h25 : T219;
  assign T219 = T289 ? 6'h24 : T220;
  assign T220 = T288 ? 6'h23 : T221;
  assign T221 = T287 ? 6'h22 : T222;
  assign T222 = T286 ? 6'h21 : T223;
  assign T223 = T285 ? 6'h20 : T224;
  assign T224 = T284 ? 5'h1f : T225;
  assign T225 = T283 ? 5'h1e : T226;
  assign T226 = T282 ? 5'h1d : T227;
  assign T227 = T281 ? 5'h1c : T228;
  assign T228 = T280 ? 5'h1b : T229;
  assign T229 = T279 ? 5'h1a : T230;
  assign T230 = T278 ? 5'h19 : T231;
  assign T231 = T277 ? 5'h18 : T232;
  assign T232 = T276 ? 5'h17 : T233;
  assign T233 = T275 ? 5'h16 : T234;
  assign T234 = T274 ? 5'h15 : T235;
  assign T235 = T273 ? 5'h14 : T236;
  assign T236 = T272 ? 5'h13 : T237;
  assign T237 = T271 ? 5'h12 : T238;
  assign T238 = T270 ? 5'h11 : T239;
  assign T239 = T269 ? 5'h10 : T240;
  assign T240 = T268 ? 4'hf : T241;
  assign T241 = T267 ? 4'he : T242;
  assign T242 = T266 ? 4'hd : T243;
  assign T243 = T265 ? 4'hc : T244;
  assign T244 = T264 ? 4'hb : T245;
  assign T245 = T263 ? 4'ha : T246;
  assign T246 = T262 ? 4'h9 : T247;
  assign T247 = T261 ? 4'h8 : T248;
  assign T248 = T260 ? 3'h7 : T249;
  assign T249 = T259 ? 3'h6 : T250;
  assign T250 = T258 ? 3'h5 : T251;
  assign T251 = T257 ? 3'h4 : T252;
  assign T252 = T256 ? 2'h3 : T253;
  assign T253 = T255 ? 2'h2 : T254;
  assign T254 = T75[1'h1];
  assign T75 = T76;
  assign T76 = remainder[6'h3f:1'h0];
  assign T255 = T75[2'h2];
  assign T256 = T75[2'h3];
  assign T257 = T75[3'h4];
  assign T258 = T75[3'h5];
  assign T259 = T75[3'h6];
  assign T260 = T75[3'h7];
  assign T261 = T75[4'h8];
  assign T262 = T75[4'h9];
  assign T263 = T75[4'ha];
  assign T264 = T75[4'hb];
  assign T265 = T75[4'hc];
  assign T266 = T75[4'hd];
  assign T267 = T75[4'he];
  assign T268 = T75[4'hf];
  assign T269 = T75[5'h10];
  assign T270 = T75[5'h11];
  assign T271 = T75[5'h12];
  assign T272 = T75[5'h13];
  assign T273 = T75[5'h14];
  assign T274 = T75[5'h15];
  assign T275 = T75[5'h16];
  assign T276 = T75[5'h17];
  assign T277 = T75[5'h18];
  assign T278 = T75[5'h19];
  assign T279 = T75[5'h1a];
  assign T280 = T75[5'h1b];
  assign T281 = T75[5'h1c];
  assign T282 = T75[5'h1d];
  assign T283 = T75[5'h1e];
  assign T284 = T75[5'h1f];
  assign T285 = T75[6'h20];
  assign T286 = T75[6'h21];
  assign T287 = T75[6'h22];
  assign T288 = T75[6'h23];
  assign T289 = T75[6'h24];
  assign T290 = T75[6'h25];
  assign T291 = T75[6'h26];
  assign T292 = T75[6'h27];
  assign T293 = T75[6'h28];
  assign T294 = T75[6'h29];
  assign T295 = T75[6'h2a];
  assign T296 = T75[6'h2b];
  assign T297 = T75[6'h2c];
  assign T298 = T75[6'h2d];
  assign T299 = T75[6'h2e];
  assign T300 = T75[6'h2f];
  assign T301 = T75[6'h30];
  assign T302 = T75[6'h31];
  assign T303 = T75[6'h32];
  assign T304 = T75[6'h33];
  assign T305 = T75[6'h34];
  assign T306 = T75[6'h35];
  assign T307 = T75[6'h36];
  assign T308 = T75[6'h37];
  assign T309 = T75[6'h38];
  assign T310 = T75[6'h39];
  assign T311 = T75[6'h3a];
  assign T312 = T75[6'h3b];
  assign T313 = T75[6'h3c];
  assign T314 = T75[6'h3d];
  assign T315 = T75[6'h3e];
  assign T316 = T75[6'h3f];
  assign T77 = 6'h3f + T317;
  assign T317 = T441 ? 6'h3f : T318;
  assign T318 = T440 ? 6'h3e : T319;
  assign T319 = T439 ? 6'h3d : T320;
  assign T320 = T438 ? 6'h3c : T321;
  assign T321 = T437 ? 6'h3b : T322;
  assign T322 = T436 ? 6'h3a : T323;
  assign T323 = T435 ? 6'h39 : T324;
  assign T324 = T434 ? 6'h38 : T325;
  assign T325 = T433 ? 6'h37 : T326;
  assign T326 = T432 ? 6'h36 : T327;
  assign T327 = T431 ? 6'h35 : T328;
  assign T328 = T430 ? 6'h34 : T329;
  assign T329 = T429 ? 6'h33 : T330;
  assign T330 = T428 ? 6'h32 : T331;
  assign T331 = T427 ? 6'h31 : T332;
  assign T332 = T426 ? 6'h30 : T333;
  assign T333 = T425 ? 6'h2f : T334;
  assign T334 = T424 ? 6'h2e : T335;
  assign T335 = T423 ? 6'h2d : T336;
  assign T336 = T422 ? 6'h2c : T337;
  assign T337 = T421 ? 6'h2b : T338;
  assign T338 = T420 ? 6'h2a : T339;
  assign T339 = T419 ? 6'h29 : T340;
  assign T340 = T418 ? 6'h28 : T341;
  assign T341 = T417 ? 6'h27 : T342;
  assign T342 = T416 ? 6'h26 : T343;
  assign T343 = T415 ? 6'h25 : T344;
  assign T344 = T414 ? 6'h24 : T345;
  assign T345 = T413 ? 6'h23 : T346;
  assign T346 = T412 ? 6'h22 : T347;
  assign T347 = T411 ? 6'h21 : T348;
  assign T348 = T410 ? 6'h20 : T349;
  assign T349 = T409 ? 5'h1f : T350;
  assign T350 = T408 ? 5'h1e : T351;
  assign T351 = T407 ? 5'h1d : T352;
  assign T352 = T406 ? 5'h1c : T353;
  assign T353 = T405 ? 5'h1b : T354;
  assign T354 = T404 ? 5'h1a : T355;
  assign T355 = T403 ? 5'h19 : T356;
  assign T356 = T402 ? 5'h18 : T357;
  assign T357 = T401 ? 5'h17 : T358;
  assign T358 = T400 ? 5'h16 : T359;
  assign T359 = T399 ? 5'h15 : T360;
  assign T360 = T398 ? 5'h14 : T361;
  assign T361 = T397 ? 5'h13 : T362;
  assign T362 = T396 ? 5'h12 : T363;
  assign T363 = T395 ? 5'h11 : T364;
  assign T364 = T394 ? 5'h10 : T365;
  assign T365 = T393 ? 4'hf : T366;
  assign T366 = T392 ? 4'he : T367;
  assign T367 = T391 ? 4'hd : T368;
  assign T368 = T390 ? 4'hc : T369;
  assign T369 = T389 ? 4'hb : T370;
  assign T370 = T388 ? 4'ha : T371;
  assign T371 = T387 ? 4'h9 : T372;
  assign T372 = T386 ? 4'h8 : T373;
  assign T373 = T385 ? 3'h7 : T374;
  assign T374 = T384 ? 3'h6 : T375;
  assign T375 = T383 ? 3'h5 : T376;
  assign T376 = T382 ? 3'h4 : T377;
  assign T377 = T381 ? 2'h3 : T378;
  assign T378 = T380 ? 2'h2 : T379;
  assign T379 = T79[1'h1];
  assign T79 = T80;
  assign T80 = divisor[6'h3f:1'h0];
  assign T380 = T79[2'h2];
  assign T381 = T79[2'h3];
  assign T382 = T79[3'h4];
  assign T383 = T79[3'h5];
  assign T384 = T79[3'h6];
  assign T385 = T79[3'h7];
  assign T386 = T79[4'h8];
  assign T387 = T79[4'h9];
  assign T388 = T79[4'ha];
  assign T389 = T79[4'hb];
  assign T390 = T79[4'hc];
  assign T391 = T79[4'hd];
  assign T392 = T79[4'he];
  assign T393 = T79[4'hf];
  assign T394 = T79[5'h10];
  assign T395 = T79[5'h11];
  assign T396 = T79[5'h12];
  assign T397 = T79[5'h13];
  assign T398 = T79[5'h14];
  assign T399 = T79[5'h15];
  assign T400 = T79[5'h16];
  assign T401 = T79[5'h17];
  assign T402 = T79[5'h18];
  assign T403 = T79[5'h19];
  assign T404 = T79[5'h1a];
  assign T405 = T79[5'h1b];
  assign T406 = T79[5'h1c];
  assign T407 = T79[5'h1d];
  assign T408 = T79[5'h1e];
  assign T409 = T79[5'h1f];
  assign T410 = T79[6'h20];
  assign T411 = T79[6'h21];
  assign T412 = T79[6'h22];
  assign T413 = T79[6'h23];
  assign T414 = T79[6'h24];
  assign T415 = T79[6'h25];
  assign T416 = T79[6'h26];
  assign T417 = T79[6'h27];
  assign T418 = T79[6'h28];
  assign T419 = T79[6'h29];
  assign T420 = T79[6'h2a];
  assign T421 = T79[6'h2b];
  assign T422 = T79[6'h2c];
  assign T423 = T79[6'h2d];
  assign T424 = T79[6'h2e];
  assign T425 = T79[6'h2f];
  assign T426 = T79[6'h30];
  assign T427 = T79[6'h31];
  assign T428 = T79[6'h32];
  assign T429 = T79[6'h33];
  assign T430 = T79[6'h34];
  assign T431 = T79[6'h35];
  assign T432 = T79[6'h36];
  assign T433 = T79[6'h37];
  assign T434 = T79[6'h38];
  assign T435 = T79[6'h39];
  assign T436 = T79[6'h3a];
  assign T437 = T79[6'h3b];
  assign T438 = T79[6'h3c];
  assign T439 = T79[6'h3d];
  assign T440 = T79[6'h3e];
  assign T441 = T79[6'h3f];
  assign T81 = T192 < T317;
  assign T82 = T94 & T83;
  assign T83 = cmdHi ? lhs_sign : T84;
  assign T84 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T85;
  assign T85 = T88 ? T87 : T86;
  assign T86 = io_req_bits_in1[5'h1f];
  assign T87 = io_req_bits_in1[6'h3f];
  assign T88 = 1'h1 == T89;
  assign T89 = io_req_bits_dw & 1'h1;
  assign lhsSigned = T90;
  assign T90 = T93 | T91;
  assign T91 = T92 == 4'h0;
  assign T92 = io_req_bits_fn & 4'h3;
  assign T93 = T61 | T17;
  assign T94 = cmdMul ^ 1'h1;
  assign T95 = isHi ? 3'h3 : 3'h5;
  assign T96 = T153 & T97;
  assign T97 = T99 | T98;
  assign T98 = count == 7'h7;
  assign T99 = T111 & T100;
  assign T100 = T101 == 64'h0;
  assign T101 = T107 & T102;
  assign T102 = ~ T103;
  assign T103 = T104[6'h3f:1'h0];
  assign T104 = $signed(65'h10000000000000000) >>> T105;
  assign T105 = T106[3'h5:1'h0];
  assign T106 = count * 4'h8;
  assign T107 = T108[6'h3f:1'h0];
  assign T108 = {T110, T109};
  assign T109 = remainder[6'h3f:1'h0];
  assign T110 = remainder[8'h81:7'h41];
  assign T111 = T113 & T112;
  assign T112 = isHi ^ 1'h1;
  assign T113 = T115 & T114;
  assign T114 = count != 7'h0;
  assign T115 = count != 7'h7;
  assign T116 = isHi ? 3'h3 : T117;
  assign T117 = neg_out ? 3'h4 : 3'h5;
  assign T118 = T162 & T119;
  assign T119 = count == 7'h40;
  assign T120 = T121 | io_kill;
  assign T121 = io_resp_ready & io_resp_valid;
  assign T122 = T123 ? 3'h1 : 3'h2;
  assign T123 = lhs_sign | T124;
  assign T124 = rhs_sign & T125;
  assign T125 = cmdMul ^ 1'h1;
  assign T442 = {66'h0, negated_remainder};
  assign T127 = state == 3'h4;
  assign T443 = {66'h0, T128};
  assign T128 = remainder[8'h80:7'h41];
  assign T129 = state == 3'h3;
  assign T130 = {T152, T131};
  assign T131 = {1'h0, T132};
  assign T132 = T133[6'h3f:1'h0];
  assign T133 = {T151, T134};
  assign T134 = T135[6'h3f:1'h0];
  assign T135 = T99 ? T147 : T136;
  assign T136 = T137;
  assign T137 = {T139, T138};
  assign T138 = T107[6'h3f:4'h8];
  assign T139 = T142 + T444;
  assign T444 = {T445, T140};
  assign T140 = T141;
  assign T141 = T108[8'h80:7'h40];
  assign T445 = T446 ? 8'hff : 8'h0;
  assign T446 = T140[7'h40];
  assign T142 = $signed(T146) * $signed(T143);
  assign T143 = T144;
  assign T144 = {1'h0, T145};
  assign T145 = T107[3'h7:1'h0];
  assign T146 = divisor;
  assign T147 = T108 >> T148;
  assign T148 = T149[3'h5:1'h0];
  assign T149 = 11'h40 - T150;
  assign T150 = count * 4'h8;
  assign T151 = T136[8'h80:7'h40];
  assign T152 = T133 >> 7'h40;
  assign T153 = T154 & isMul;
  assign T154 = state == 3'h2;
  assign T447 = {1'h0, T155};
  assign T155 = {T159, T156};
  assign T156 = {T158, T157};
  assign T157 = less ^ 1'h1;
  assign T158 = remainder[6'h3f:1'h0];
  assign T159 = less ? T161 : T160;
  assign T160 = subtractor[6'h3f:1'h0];
  assign T161 = remainder[7'h7f:7'h40];
  assign T162 = T164 & T163;
  assign T163 = isMul ^ 1'h1;
  assign T164 = state == 3'h2;
  assign T448 = {3'h0, T165};
  assign T165 = T166 << T71;
  assign T166 = remainder[6'h3f:1'h0];
  assign T167 = T162 & T168;
  assign T168 = T171 & T169;
  assign T169 = T170 | T81;
  assign T170 = 6'h0 < T73;
  assign T171 = T172 & less;
  assign T172 = count == 7'h0;
  assign T449 = {66'h0, lhs_in};
  assign lhs_in = {T174, T173};
  assign T173 = io_req_bits_in1[5'h1f:1'h0];
  assign T174 = T177 ? T176 : T175;
  assign T175 = 32'h0 - T450;
  assign T450 = {31'h0, lhs_sign};
  assign T176 = io_req_bits_in1[6'h3f:6'h20];
  assign T177 = 1'h1 == T178;
  assign T178 = io_req_bits_dw & 1'h1;
  assign T179 = {T181, T180};
  assign T180 = remainder[5'h1f:1'h0];
  assign T181 = 32'h0 - T451;
  assign T451 = {31'h0, T182};
  assign T182 = remainder[5'h1f];
  assign T183 = 1'h0 == T184;
  assign T184 = req_dw & 1'h1;
  assign T185 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T186;
  assign T186 = state == 3'h5;
  assign io_req_ready = T187;
  assign T187 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T449;
    end else if(T167) begin
      remainder <= T448;
    end else if(T162) begin
      remainder <= T447;
    end else if(T153) begin
      remainder <= T130;
    end else if(T129) begin
      remainder <= T443;
    end else if(T127) begin
      remainder <= T442;
    end else if(T11) begin
      remainder <= T188;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T122;
    end else if(T120) begin
      state <= 3'h0;
    end else if(T118) begin
      state <= T116;
    end else if(T96) begin
      state <= T95;
    end else if(T129) begin
      state <= T28;
    end else if(T127) begin
      state <= 3'h5;
    end else if(T20) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T82;
    end else if(T31) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T48;
    end else if(T45) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T167) begin
      count <= T191;
    end else if(T162) begin
      count <= T70;
    end else if(T153) begin
      count <= T69;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module Rocket(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    output io_imem_req_valid,
    output[39:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [39:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [38:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_btb_update_bits_pc,
    output[38:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output[38:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_bht_update_bits_prediction_bits_target,
    output[5:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output[38:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_ras_update_bits_prediction_bits_target,
    output[5:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    output io_imem_invalidate,
    input [39:0] io_imem_npc,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output[39:0] io_dmem_req_bits_addr,
    output[9:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_kill,
    output io_dmem_req_bits_phys,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [39:0] io_dmem_resp_bits_addr,
    input [9:0] io_dmem_resp_bits_tag,
    input [4:0] io_dmem_resp_bits_cmd,
    input [2:0] io_dmem_resp_bits_typ,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_word_bypass,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [9:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    output io_dmem_invalidate_lr,
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_status_sd,
    output[30:0] io_ptw_status_zero2,
    output io_ptw_status_sd_rv32,
    output[8:0] io_ptw_status_zero1,
    output[4:0] io_ptw_status_vm,
    output io_ptw_status_mprv,
    output[1:0] io_ptw_status_xs,
    output[1:0] io_ptw_status_fs,
    output[1:0] io_ptw_status_prv3,
    output io_ptw_status_ie3,
    output[1:0] io_ptw_status_prv2,
    output io_ptw_status_ie2,
    output[1:0] io_ptw_status_prv1,
    output io_ptw_status_ie1,
    output[1:0] io_ptw_status_prv,
    output io_ptw_status_ie,
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    output io_fpu_valid,
    input  io_fpu_fcsr_rdy,
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input  io_fpu_dec_ldst,
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    input  io_fpu_dec_swap12,
    input  io_fpu_dec_swap23,
    input  io_fpu_dec_single,
    input  io_fpu_dec_fromint,
    input  io_fpu_dec_toint,
    input  io_fpu_dec_fastpipe,
    input  io_fpu_dec_fma,
    input  io_fpu_dec_div,
    input  io_fpu_dec_sqrt,
    input  io_fpu_dec_round,
    input  io_fpu_dec_wflags,
    input  io_fpu_sboard_set,
    input  io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input  io_fpu_cp_req_ready,
    //output io_fpu_cp_req_valid
    //output[4:0] io_fpu_cp_req_bits_cmd
    //output io_fpu_cp_req_bits_ldst
    //output io_fpu_cp_req_bits_wen
    //output io_fpu_cp_req_bits_ren1
    //output io_fpu_cp_req_bits_ren2
    //output io_fpu_cp_req_bits_ren3
    //output io_fpu_cp_req_bits_swap12
    //output io_fpu_cp_req_bits_swap23
    //output io_fpu_cp_req_bits_single
    //output io_fpu_cp_req_bits_fromint
    //output io_fpu_cp_req_bits_toint
    //output io_fpu_cp_req_bits_fastpipe
    //output io_fpu_cp_req_bits_fma
    //output io_fpu_cp_req_bits_div
    //output io_fpu_cp_req_bits_sqrt
    //output io_fpu_cp_req_bits_round
    //output io_fpu_cp_req_bits_wflags
    //output[2:0] io_fpu_cp_req_bits_rm
    //output[1:0] io_fpu_cp_req_bits_typ
    //output[64:0] io_fpu_cp_req_bits_in1
    //output[64:0] io_fpu_cp_req_bits_in2
    //output[64:0] io_fpu_cp_req_bits_in3
    //output io_fpu_cp_resp_ready
    input  io_fpu_cp_resp_valid,
    input [64:0] io_fpu_cp_resp_bits_data,
    //input [4:0] io_fpu_cp_resp_bits_exc
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    output io_rocc_resp_ready,
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [9:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[9:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[9:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_autl_acquire_ready
    input  io_rocc_autl_acquire_valid,
    input [25:0] io_rocc_autl_acquire_bits_addr_block,
    input [5:0] io_rocc_autl_acquire_bits_client_xact_id,
    input [1:0] io_rocc_autl_acquire_bits_addr_beat,
    input  io_rocc_autl_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_autl_acquire_bits_a_type,
    input [16:0] io_rocc_autl_acquire_bits_union,
    input [127:0] io_rocc_autl_acquire_bits_data,
    input  io_rocc_autl_grant_ready,
    //output io_rocc_autl_grant_valid
    //output[1:0] io_rocc_autl_grant_bits_addr_beat
    //output[5:0] io_rocc_autl_grant_bits_client_xact_id
    //output[3:0] io_rocc_autl_grant_bits_manager_xact_id
    //output io_rocc_autl_grant_bits_is_builtin_type
    //output[3:0] io_rocc_autl_grant_bits_g_type
    //output[127:0] io_rocc_autl_grant_bits_data
    //output io_rocc_fpu_req_ready
    input  io_rocc_fpu_req_valid,
    input [4:0] io_rocc_fpu_req_bits_cmd,
    input  io_rocc_fpu_req_bits_ldst,
    input  io_rocc_fpu_req_bits_wen,
    input  io_rocc_fpu_req_bits_ren1,
    input  io_rocc_fpu_req_bits_ren2,
    input  io_rocc_fpu_req_bits_ren3,
    input  io_rocc_fpu_req_bits_swap12,
    input  io_rocc_fpu_req_bits_swap23,
    input  io_rocc_fpu_req_bits_single,
    input  io_rocc_fpu_req_bits_fromint,
    input  io_rocc_fpu_req_bits_toint,
    input  io_rocc_fpu_req_bits_fastpipe,
    input  io_rocc_fpu_req_bits_fma,
    input  io_rocc_fpu_req_bits_div,
    input  io_rocc_fpu_req_bits_sqrt,
    input  io_rocc_fpu_req_bits_round,
    input  io_rocc_fpu_req_bits_wflags,
    input [2:0] io_rocc_fpu_req_bits_rm,
    input [1:0] io_rocc_fpu_req_bits_typ,
    input [64:0] io_rocc_fpu_req_bits_in1,
    input [64:0] io_rocc_fpu_req_bits_in2,
    input [64:0] io_rocc_fpu_req_bits_in3,
    input  io_rocc_fpu_resp_ready,
    //output io_rocc_fpu_resp_valid
    //output[64:0] io_rocc_fpu_resp_bits_data
    //output[4:0] io_rocc_fpu_resp_bits_exc
    output io_rocc_exception,
    output[11:0] io_rocc_csr_waddr,
    output[63:0] io_rocc_csr_wdata,
    output io_rocc_csr_wen
    //output io_rocc_host_id
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  wire ctrl_killd;
  wire T7;
  wire T8;
  wire ctrl_stalld;
  wire T9;
  wire id_do_fence;
  wire T10;
  wire T11;
  wire id_csr_en;
  wire[2:0] id_ctrl_csr;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire[31:0] T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire[31:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire id_ctrl_rocc;
  wire T23;
  wire T24;
  wire[31:0] T25;
  wire T26;
  wire[31:0] T27;
  wire id_ctrl_mem;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire T41;
  wire[31:0] T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  reg  id_reg_fence;
  wire T1072;
  wire T48;
  wire T49;
  wire id_fence_next;
  wire T50;
  wire id_amo_rl;
  wire id_ctrl_amo;
  wire T51;
  wire[31:0] T52;
  wire id_ctrl_fence;
  wire T53;
  wire[31:0] T54;
  wire T55;
  wire id_ctrl_fence_i;
  wire T56;
  wire[31:0] T57;
  wire T58;
  wire id_amo_aq;
  wire id_mem_busy;
  wire T59;
  wire T60;
  wire id_rocc_busy;
  wire T61;
  reg  wb_ctrl_rocc;
  wire T62;
  reg  mem_ctrl_rocc;
  wire T63;
  reg  ex_ctrl_rocc;
  wire T64;
  wire T65;
  reg  wb_reg_valid;
  wire T66;
  wire ctrl_killm;
  wire fpu_kill_mem;
  wire T67;
  reg  mem_ctrl_fp;
  wire T68;
  reg  ex_ctrl_fp;
  wire T69;
  wire id_ctrl_fp;
  wire T70;
  wire T71;
  wire[31:0] T72;
  wire T73;
  wire T74;
  wire[31:0] T75;
  wire T76;
  wire[31:0] T77;
  reg  mem_reg_valid;
  wire T78;
  wire ctrl_killx;
  wire T79;
  reg  ex_reg_valid;
  wire T80;
  wire T81;
  wire replay_ex;
  wire T82;
  wire replay_ex_load_use;
  reg  ex_reg_load_use;
  wire T83;
  wire id_load_use;
  wire T84;
  reg  mem_ctrl_mem;
  wire T85;
  reg  ex_ctrl_mem;
  wire T86;
  wire T87;
  wire data_hazard_mem;
  wire T88;
  wire T89;
  wire T90;
  wire[4:0] mem_waddr;
  wire[4:0] id_waddr;
  wire T91;
  wire T92;
  wire id_ctrl_wxd;
  wire T93;
  wire T94;
  wire[31:0] T95;
  wire T96;
  wire T97;
  wire[31:0] T98;
  wire T99;
  wire T100;
  wire[31:0] T101;
  wire T102;
  wire T103;
  wire[31:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[31:0] T108;
  wire T109;
  wire T110;
  wire[31:0] T111;
  wire T112;
  wire T113;
  wire[31:0] T114;
  wire T115;
  wire T116;
  wire[31:0] T117;
  wire T118;
  wire[31:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[4:0] id_raddr_1;
  wire T123;
  wire T124;
  wire id_ctrl_rxs2;
  wire T125;
  wire T126;
  wire[31:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire T133;
  wire[31:0] T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire T138;
  wire[4:0] id_raddr_0;
  wire T139;
  wire T140;
  wire id_ctrl_rxs1;
  wire T141;
  wire T142;
  wire[31:0] T143;
  wire T144;
  wire T145;
  wire[31:0] T146;
  wire T147;
  wire T148;
  wire[31:0] T149;
  wire T150;
  wire T151;
  wire[31:0] T152;
  wire T153;
  wire T154;
  wire[31:0] T155;
  wire T156;
  wire T157;
  wire[31:0] T158;
  wire T159;
  wire[31:0] T160;
  reg  mem_ctrl_wxd;
  wire T161;
  reg  ex_ctrl_wxd;
  wire T162;
  wire wb_dcache_miss;
  wire T163;
  reg  wb_ctrl_mem;
  wire T164;
  wire replay_ex_structural;
  wire T165;
  wire T166;
  reg  ex_ctrl_div;
  wire T167;
  wire id_ctrl_div;
  wire T168;
  wire[31:0] T169;
  wire T170;
  wire T171;
  wire take_pc;
  wire take_pc_mem;
  wire T172;
  wire T173;
  wire mem_npc_misaligned;
  wire[39:0] mem_npc;
  wire[39:0] T174;
  wire[39:0] T175;
  wire[39:0] mem_br_target;
  wire[39:0] T1073;
  wire[21:0] T176;
  wire[21:0] T177;
  wire[21:0] T178;
  wire[21:0] T179;
  wire[11:0] T180;
  wire[4:0] T181;
  wire[3:0] T182;
  wire[6:0] T183;
  wire[5:0] T184;
  wire T185;
  wire T186;
  wire[9:0] T187;
  wire[8:0] T188;
  wire[7:0] T189;
  wire[7:0] T190;
  wire T191;
  wire T192;
  reg  mem_ctrl_jal;
  wire T193;
  reg  ex_ctrl_jal;
  wire T194;
  wire id_ctrl_jal;
  wire[21:0] T1074;
  wire[14:0] T195;
  wire[14:0] T196;
  wire[11:0] T197;
  wire[4:0] T198;
  wire[3:0] T199;
  wire[6:0] T200;
  wire[5:0] T201;
  wire T202;
  wire T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire T207;
  wire[6:0] T1075;
  wire T1076;
  wire T208;
  wire mem_br_taken;
  reg [63:0] bypass_mux_1;
  wire[63:0] T209;
  reg  mem_ctrl_branch;
  wire T210;
  reg  ex_ctrl_branch;
  wire T211;
  wire id_ctrl_branch;
  wire T212;
  wire[31:0] T213;
  wire[17:0] T1077;
  wire T1078;
  wire[39:0] T214;
  reg [39:0] mem_reg_pc;
  wire[39:0] T215;
  reg [39:0] ex_reg_pc;
  wire[39:0] T216;
  wire[39:0] T217;
  wire[39:0] T218;
  wire[38:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire[1:0] T225;
  wire T226;
  wire T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire T230;
  wire[25:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  reg  mem_ctrl_jalr;
  wire T236;
  reg  ex_ctrl_jalr;
  wire T237;
  wire id_ctrl_jalr;
  wire T238;
  wire[31:0] T239;
  wire want_take_pc_mem;
  wire T240;
  reg  mem_reg_flush_pipe;
  wire T241;
  reg  ex_reg_flush_pipe;
  wire T242;
  wire T243;
  wire id_csr_flush;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  wire[11:0] id_csr_addr;
  wire T249;
  wire T250;
  wire id_csr_ren;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire id_system_insn;
  wire mem_misprediction;
  wire T255;
  wire T256;
  wire T257;
  wire mem_wrong_npc;
  wire T258;
  wire T259;
  wire take_pc_wb;
  wire T260;
  wire T261;
  wire wb_xcpt;
  reg  wb_reg_xcpt;
  wire T262;
  wire T263;
  wire mem_xcpt;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  reg  mem_reg_xcpt;
  wire T278;
  wire ex_xcpt;
  wire T279;
  wire T280;
  reg  ex_reg_xcpt;
  wire T281;
  wire id_xcpt;
  wire id_illegal_insn;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire id_ctrl_legal;
  wire T290;
  wire T291;
  wire[31:0] T292;
  wire T293;
  wire T294;
  wire[31:0] T295;
  wire T296;
  wire T297;
  wire[31:0] T298;
  wire T299;
  wire T300;
  wire[31:0] T301;
  wire T302;
  wire T303;
  wire[31:0] T304;
  wire T305;
  wire T306;
  wire[31:0] T307;
  wire T308;
  wire T309;
  wire[31:0] T310;
  wire T311;
  wire T312;
  wire[31:0] T313;
  wire T314;
  wire T315;
  wire[31:0] T316;
  wire T317;
  wire T318;
  wire[31:0] T319;
  wire T320;
  wire T321;
  wire[31:0] T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire[31:0] T327;
  wire T328;
  wire T329;
  wire[31:0] T330;
  wire T331;
  wire T332;
  wire[31:0] T333;
  wire T334;
  wire T335;
  wire[31:0] T336;
  wire T337;
  wire T338;
  wire T339;
  wire[31:0] T340;
  wire T341;
  wire T342;
  wire T343;
  wire[31:0] T344;
  wire T345;
  wire T346;
  wire[31:0] T347;
  wire T348;
  wire T349;
  wire[31:0] T350;
  wire T351;
  wire T352;
  wire[31:0] T353;
  wire T354;
  wire T355;
  wire[31:0] T356;
  wire T357;
  wire T358;
  wire[31:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire[31:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire[31:0] T370;
  wire T371;
  wire T372;
  wire[31:0] T373;
  wire T374;
  wire T375;
  wire[31:0] T376;
  wire T377;
  wire T378;
  wire[31:0] T379;
  wire T380;
  wire T381;
  wire[31:0] T382;
  wire T383;
  wire T384;
  wire[31:0] T385;
  wire T386;
  wire T387;
  wire[31:0] T388;
  wire T389;
  wire T390;
  wire[31:0] T391;
  wire T392;
  wire T393;
  wire[31:0] T394;
  wire T395;
  wire T396;
  wire[31:0] T397;
  wire T398;
  wire T399;
  wire[31:0] T400;
  wire T401;
  wire T402;
  wire[31:0] T403;
  wire T404;
  wire T405;
  wire[31:0] T406;
  wire T407;
  wire T408;
  wire[31:0] T409;
  wire T410;
  wire T411;
  reg  ex_reg_xcpt_interrupt;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  reg  mem_reg_xcpt_interrupt;
  wire T416;
  wire T417;
  wire replay_wb;
  wire T418;
  wire T419;
  wire T420;
  wire replay_wb_common;
  reg  wb_reg_replay;
  wire T421;
  wire T422;
  wire replay_mem;
  wire T423;
  reg  mem_reg_replay;
  wire T424;
  wire T425;
  wire dcache_kill_mem;
  wire T426;
  wire T427;
  wire killm_common;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  reg  wb_reg_rocc_pending;
  wire T1079;
  wire T439;
  wire T440;
  wire T441;
  wire wb_rocc_val;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire id_stall_fpu;
  wire T449;
  wire T450;
  wire T451;
  reg [31:0] R452;
  wire[31:0] T1080;
  wire[31:0] T453;
  wire[31:0] T454;
  wire[31:0] T455;
  wire[31:0] T456;
  wire[31:0] T457;
  wire[31:0] T458;
  wire[4:0] wb_waddr;
  wire T459;
  wire wb_valid;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg  wb_ctrl_wfd;
  wire T465;
  reg  mem_ctrl_wfd;
  wire T466;
  reg  ex_ctrl_wfd;
  wire T467;
  wire id_ctrl_wfd;
  wire T468;
  wire T469;
  wire[31:0] T470;
  wire T471;
  wire T472;
  wire T473;
  wire[31:0] T474;
  wire T475;
  wire[31:0] T476;
  wire[31:0] T477;
  wire[31:0] T478;
  wire[31:0] T479;
  wire[31:0] T480;
  wire[4:0] dmem_resp_waddr;
  wire[9:0] T481;
  wire T482;
  wire dmem_resp_fpu;
  wire T483;
  wire dmem_resp_replay;
  wire T484;
  wire[31:0] T485;
  wire[31:0] T486;
  wire[31:0] T487;
  wire[31:0] T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire[4:0] id_raddr3;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire id_sboard_hazard;
  wire T501;
  wire T502;
  wire[31:0] T503;
  wire[31:0] T504;
  wire[31:0] T505;
  wire[31:0] T506;
  wire[4:0] ll_waddr;
  wire[4:0] T507;
  wire[4:0] T508;
  wire T509;
  wire T510;
  wire dmem_resp_xpu;
  wire T511;
  wire T512;
  wire ll_wen;
  wire T513;
  wire T514;
  wire T515;
  reg [31:0] R516;
  wire[31:0] T1081;
  wire[31:0] T517;
  wire[31:0] T518;
  wire[31:0] T519;
  wire[31:0] T520;
  wire[31:0] T521;
  wire T522;
  wire wb_wen;
  reg  wb_ctrl_wxd;
  wire T523;
  wire wb_set_sboard;
  wire T524;
  reg  wb_ctrl_div;
  wire T525;
  reg  mem_ctrl_div;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire id_wb_hazard;
  wire T534;
  wire fp_data_hazard_wb;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire data_hazard_wb;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire id_mem_hazard;
  wire T556;
  wire fp_data_hazard_mem;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire mem_cannot_bypass;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  reg  mem_mem_cmd_bh;
  wire T573;
  wire ex_slow_bypass;
  wire T574;
  wire T575;
  reg [2:0] ex_ctrl_mem_type;
  wire[2:0] T576;
  wire[2:0] id_ctrl_mem_type;
  wire[2:0] T577;
  wire[1:0] T578;
  wire T579;
  wire[31:0] T580;
  wire T581;
  wire[31:0] T582;
  wire T583;
  wire[31:0] T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  reg [4:0] ex_ctrl_mem_cmd;
  wire[4:0] T591;
  wire[4:0] id_ctrl_mem_cmd;
  wire[4:0] T592;
  wire[3:0] T593;
  wire[2:0] T594;
  wire[1:0] T595;
  wire T596;
  wire T597;
  wire[31:0] T598;
  wire T599;
  wire T600;
  wire[31:0] T601;
  wire T602;
  wire[31:0] T603;
  wire T604;
  wire T605;
  wire[31:0] T606;
  wire T607;
  wire[31:0] T608;
  wire T609;
  wire T610;
  wire[31:0] T611;
  wire T612;
  wire T613;
  wire[31:0] T614;
  wire T615;
  wire[31:0] T616;
  wire T617;
  reg [2:0] mem_ctrl_csr;
  wire[2:0] T618;
  reg [2:0] ex_ctrl_csr;
  wire[2:0] T619;
  wire[2:0] T620;
  wire[2:0] id_csr;
  wire id_ex_hazard;
  wire T621;
  wire fp_data_hazard_ex;
  wire T622;
  wire T623;
  wire T624;
  wire[4:0] ex_waddr;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire ex_cannot_bypass;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire data_hazard_ex;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[31:0] T652;
  wire[63:0] T653;
  reg [63:0] R654;
  reg [63:0] R655;
  wire[63:0] ex_rs_1;
  wire[63:0] T656;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire[1:0] T671;
  wire[63:0] id_rs_1;
  wire[63:0] T672;
  wire[63:0] T673;
  reg [63:0] T674 [30:0];
  wire[63:0] T675;
  wire T676;
  wire T677;
  wire[4:0] T678;
  wire T679;
  wire T680;
  wire[4:0] rf_waddr;
  wire rf_wen;
  wire[4:0] T681;
  wire[4:0] T682;
  wire[4:0] T683;
  wire[63:0] rf_wdata;
  wire[63:0] T684;
  wire[63:0] T685;
  reg [63:0] bypass_mux_2;
  wire[63:0] T686;
  wire[63:0] T687;
  wire[63:0] mem_int_wdata;
  wire[63:0] T688;
  wire[63:0] T689;
  wire[63:0] T1082;
  wire[23:0] T1083;
  wire T1084;
  wire T690;
  wire T691;
  reg [2:0] wb_ctrl_csr;
  wire[2:0] T692;
  wire[63:0] ll_wdata;
  wire[63:0] T693;
  wire T694;
  wire dmem_resp_valid;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T706;
  wire[61:0] T707;
  wire[63:0] T708;
  wire[63:0] T709;
  wire T710;
  wire[1:0] T711;
  wire[63:0] T712;
  wire T713;
  wire T714;
  reg  ex_reg_rs_bypass_1;
  wire T715;
  wire[4:0] T716;
  wire[4:0] T717;
  wire[63:0] T718;
  reg [63:0] R719;
  reg [63:0] R720;
  wire[63:0] ex_rs_0;
  wire[63:0] T721;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire[1:0] T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[63:0] id_rs_0;
  wire[63:0] T733;
  wire[63:0] T734;
  wire[4:0] T735;
  wire[4:0] T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T747;
  wire[61:0] T748;
  wire[63:0] T749;
  wire[63:0] T750;
  wire T751;
  wire[1:0] T752;
  wire[63:0] T753;
  wire T754;
  wire T755;
  reg  ex_reg_rs_bypass_0;
  wire T756;
  wire[4:0] T757;
  wire[4:0] T758;
  wire T759;
  wire[63:0] T760;
  wire[4:0] T761;
  wire[4:0] T762;
  wire[39:0] T763;
  reg [39:0] wb_reg_pc;
  wire[39:0] T764;
  wire T765;
  wire[32:0] T766;
  wire[32:0] T767;
  wire T768;
  wire[1127:0] T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  reg  R775;
  wire T776;
  reg  ex_ctrl_alu_dw;
  wire T777;
  wire id_ctrl_alu_dw;
  wire T778;
  wire T779;
  wire[31:0] T780;
  wire T781;
  wire T782;
  wire[31:0] T783;
  wire T784;
  wire[31:0] T785;
  reg [3:0] ex_ctrl_alu_fn;
  wire[3:0] T786;
  wire[3:0] id_ctrl_alu_fn;
  wire[3:0] T787;
  wire[2:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire[31:0] T792;
  wire T793;
  wire T794;
  wire[31:0] T795;
  wire T796;
  wire[31:0] T797;
  wire T798;
  wire T799;
  wire[31:0] T800;
  wire T801;
  wire T802;
  wire[31:0] T803;
  wire T804;
  wire T805;
  wire[31:0] T806;
  wire T807;
  wire T808;
  wire[31:0] T809;
  wire T810;
  wire T811;
  wire[31:0] T812;
  wire T813;
  wire[31:0] T814;
  wire T815;
  wire T816;
  wire[31:0] T817;
  wire T818;
  wire T819;
  wire[31:0] T820;
  wire T821;
  wire T822;
  wire[31:0] T823;
  wire T824;
  wire[31:0] T825;
  wire T826;
  wire T827;
  wire[31:0] T828;
  wire T829;
  wire T830;
  wire T831;
  wire[31:0] T832;
  wire T833;
  wire[63:0] T834;
  wire[63:0] ex_op1;
  wire[63:0] T1085;
  wire[39:0] T835;
  wire[39:0] T836;
  wire T837;
  reg [1:0] ex_ctrl_sel_alu1;
  wire[1:0] T838;
  wire[1:0] id_ctrl_sel_alu1;
  wire[1:0] T839;
  wire T840;
  wire T841;
  wire[31:0] T842;
  wire T843;
  wire T844;
  wire[31:0] T845;
  wire T846;
  wire T847;
  wire[31:0] T848;
  wire T849;
  wire T850;
  wire[31:0] T851;
  wire T852;
  wire T853;
  wire[31:0] T854;
  wire T855;
  wire[31:0] T856;
  wire T857;
  wire T858;
  wire[31:0] T859;
  wire T860;
  wire[31:0] T861;
  wire[23:0] T1086;
  wire T1087;
  wire[63:0] T862;
  wire T863;
  wire[63:0] T864;
  wire[63:0] ex_op2;
  wire[63:0] T1088;
  wire[31:0] T865;
  wire[31:0] T1089;
  wire[3:0] T866;
  wire T867;
  reg [1:0] ex_ctrl_sel_alu2;
  wire[1:0] T868;
  wire[1:0] id_ctrl_sel_alu2;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire[31:0] T872;
  wire T873;
  wire T874;
  wire T875;
  wire[31:0] T876;
  wire T877;
  wire T878;
  wire[31:0] T879;
  wire T880;
  wire T881;
  wire[31:0] T882;
  wire T883;
  wire[27:0] T1090;
  wire T1091;
  wire[31:0] ex_imm;
  wire[31:0] T884;
  wire[11:0] T885;
  wire[4:0] T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  reg [2:0] ex_ctrl_sel_imm;
  wire[2:0] T892;
  wire[2:0] id_ctrl_sel_imm;
  wire[2:0] T893;
  wire[1:0] T894;
  wire T895;
  wire T896;
  wire[31:0] T897;
  wire T898;
  wire[31:0] T899;
  wire T900;
  wire T901;
  wire[31:0] T902;
  wire T903;
  wire T904;
  wire[31:0] T905;
  wire T906;
  wire T907;
  wire[31:0] T908;
  wire T909;
  wire[31:0] T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[3:0] T918;
  wire[3:0] T919;
  wire T920;
  wire[3:0] T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire[6:0] T926;
  wire[5:0] T927;
  wire[5:0] T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[19:0] T948;
  wire[18:0] T949;
  wire[7:0] T950;
  wire[7:0] T951;
  wire[7:0] T952;
  wire[7:0] T1092;
  wire T953;
  wire T954;
  wire T955;
  wire[10:0] T956;
  wire[10:0] T1093;
  wire[10:0] T957;
  wire[10:0] T958;
  wire T959;
  wire T960;
  wire[31:0] T1094;
  wire T1095;
  wire[63:0] T961;
  wire T962;
  reg [63:0] wb_reg_cause;
  wire[63:0] T963;
  wire[63:0] mem_cause;
  wire[63:0] T1096;
  wire[2:0] T964;
  wire[2:0] T965;
  wire[2:0] T966;
  wire[2:0] T967;
  reg [63:0] mem_reg_cause;
  wire[63:0] T968;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T969;
  wire[63:0] id_cause;
  wire[63:0] T1097;
  wire[1:0] T970;
  wire[2:0] T971;
  wire[11:0] T972;
  wire T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T979;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T980;
  wire T981;
  wire T982;
  wire T983;
  reg  ex_ctrl_rxs2;
  wire T984;
  wire T985;
  wire[6:0] T986;
  wire[4:0] T987;
  wire T988;
  wire T989;
  wire T990;
  wire[4:0] T991;
  wire[4:0] T992;
  wire[6:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire[63:0] T997;
  wire T998;
  wire[9:0] T1098;
  wire[5:0] T999;
  wire[39:0] T1000;
  wire[39:0] T1001;
  wire[38:0] T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire[1:0] T1006;
  wire T1007;
  wire[1:0] T1008;
  wire T1009;
  wire T1010;
  wire[25:0] T1011;
  wire[25:0] T1012;
  wire T1013;
  wire[25:0] T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  reg  wb_ctrl_fence_i;
  wire T1021;
  reg  mem_ctrl_fence_i;
  wire T1022;
  reg  ex_ctrl_fence_i;
  wire T1023;
  wire[38:0] T1099;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire[38:0] T1100;
  wire T1031;
  wire T1032;
  wire T1033;
  wire[38:0] T1101;
  wire T1034;
  wire T1035;
  wire[4:0] T1036;
  wire[4:0] T1037;
  wire T1038;
  wire[38:0] T1102;
  wire[38:0] T1103;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T1039;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T1040;
  wire T1041;
  wire T1042;
  reg  ex_reg_btb_hit;
  wire T1043;
  reg [6:0] mem_reg_btb_resp_bht_history;
  wire[6:0] T1044;
  reg [6:0] ex_reg_btb_resp_bht_history;
  wire[6:0] T1045;
  reg [5:0] mem_reg_btb_resp_entry;
  wire[5:0] T1046;
  reg [5:0] ex_reg_btb_resp_entry;
  wire[5:0] T1047;
  reg [38:0] mem_reg_btb_resp_target;
  wire[38:0] T1048;
  reg [38:0] ex_reg_btb_resp_target;
  wire[38:0] T1049;
  reg  mem_reg_btb_resp_bridx;
  wire T1050;
  reg  ex_reg_btb_resp_bridx;
  wire T1051;
  reg  mem_reg_btb_resp_mask;
  wire T1052;
  reg  ex_reg_btb_resp_mask;
  wire T1053;
  reg  mem_reg_btb_resp_taken;
  wire T1054;
  reg  ex_reg_btb_resp_taken;
  wire T1055;
  reg  mem_reg_btb_hit;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[39:0] T1068;
  wire[39:0] T1069;
  wire[39:0] T1070;
  wire T1071;
  wire csr_io_host_csr_req_ready;
  wire csr_io_host_csr_resp_valid;
  wire[63:0] csr_io_host_csr_resp_bits;
  wire csr_io_host_debug_stats_csr;
  wire[63:0] csr_io_rw_rdata;
  wire csr_io_csr_stall;
  wire csr_io_csr_xcpt;
  wire csr_io_eret;
  wire csr_io_status_sd;
  wire[30:0] csr_io_status_zero2;
  wire csr_io_status_sd_rv32;
  wire[8:0] csr_io_status_zero1;
  wire[4:0] csr_io_status_vm;
  wire csr_io_status_mprv;
  wire[1:0] csr_io_status_xs;
  wire[1:0] csr_io_status_fs;
  wire[1:0] csr_io_status_prv3;
  wire csr_io_status_ie3;
  wire[1:0] csr_io_status_prv2;
  wire csr_io_status_ie2;
  wire[1:0] csr_io_status_prv1;
  wire csr_io_status_ie1;
  wire[1:0] csr_io_status_prv;
  wire csr_io_status_ie;
  wire[31:0] csr_io_ptbr;
  wire[39:0] csr_io_evec;
  wire csr_io_fatc;
  wire[63:0] csr_io_time;
  wire[2:0] csr_io_fcsr_rm;
  wire[11:0] csr_io_rocc_csr_waddr;
  wire[63:0] csr_io_rocc_csr_wdata;
  wire csr_io_rocc_csr_wen;
  wire csr_io_interrupt;
  wire[63:0] csr_io_interrupt_cause;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    id_reg_fence = {1{$random}};
    wb_ctrl_rocc = {1{$random}};
    mem_ctrl_rocc = {1{$random}};
    ex_ctrl_rocc = {1{$random}};
    wb_reg_valid = {1{$random}};
    mem_ctrl_fp = {1{$random}};
    ex_ctrl_fp = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_ctrl_mem = {1{$random}};
    ex_ctrl_mem = {1{$random}};
    mem_ctrl_wxd = {1{$random}};
    ex_ctrl_wxd = {1{$random}};
    wb_ctrl_mem = {1{$random}};
    ex_ctrl_div = {1{$random}};
    mem_ctrl_jal = {1{$random}};
    ex_ctrl_jal = {1{$random}};
    bypass_mux_1 = {2{$random}};
    mem_ctrl_branch = {1{$random}};
    ex_ctrl_branch = {1{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    mem_ctrl_jalr = {1{$random}};
    ex_ctrl_jalr = {1{$random}};
    mem_reg_flush_pipe = {1{$random}};
    ex_reg_flush_pipe = {1{$random}};
    wb_reg_xcpt = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    wb_reg_replay = {1{$random}};
    mem_reg_replay = {1{$random}};
    wb_reg_rocc_pending = {1{$random}};
    R452 = {1{$random}};
    wb_ctrl_wfd = {1{$random}};
    mem_ctrl_wfd = {1{$random}};
    ex_ctrl_wfd = {1{$random}};
    R516 = {1{$random}};
    wb_ctrl_wxd = {1{$random}};
    wb_ctrl_div = {1{$random}};
    mem_ctrl_div = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_ctrl_mem_type = {1{$random}};
    ex_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_csr = {1{$random}};
    ex_ctrl_csr = {1{$random}};
    R654 = {2{$random}};
    R655 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T674[initvar] = {2{$random}};
    bypass_mux_2 = {2{$random}};
    wb_ctrl_csr = {1{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R719 = {2{$random}};
    R720 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    R775 = {1{$random}};
    ex_ctrl_alu_dw = {1{$random}};
    ex_ctrl_alu_fn = {1{$random}};
    ex_ctrl_sel_alu1 = {1{$random}};
    ex_ctrl_sel_alu2 = {1{$random}};
    ex_ctrl_sel_imm = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
    ex_ctrl_rxs2 = {1{$random}};
    wb_ctrl_fence_i = {1{$random}};
    mem_ctrl_fence_i = {1{$random}};
    ex_ctrl_fence_i = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_bridx = {1{$random}};
    ex_reg_btb_resp_bridx = {1{$random}};
    mem_reg_btb_resp_mask = {1{$random}};
    ex_reg_btb_resp_mask = {1{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_host_id = {1{$random}};
//  assign io_rocc_fpu_resp_bits_exc = {1{$random}};
//  assign io_rocc_fpu_resp_bits_data = {3{$random}};
//  assign io_rocc_fpu_resp_valid = {1{$random}};
//  assign io_rocc_fpu_req_ready = {1{$random}};
//  assign io_rocc_autl_grant_bits_data = {4{$random}};
//  assign io_rocc_autl_grant_bits_g_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_autl_grant_valid = {1{$random}};
//  assign io_rocc_autl_acquire_ready = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_fpu_cp_resp_ready = {1{$random}};
//  assign io_fpu_cp_req_bits_in3 = {3{$random}};
//  assign io_fpu_cp_req_bits_in2 = {3{$random}};
//  assign io_fpu_cp_req_bits_in1 = {3{$random}};
//  assign io_fpu_cp_req_bits_typ = {1{$random}};
//  assign io_fpu_cp_req_bits_rm = {1{$random}};
//  assign io_fpu_cp_req_bits_wflags = {1{$random}};
//  assign io_fpu_cp_req_bits_round = {1{$random}};
//  assign io_fpu_cp_req_bits_sqrt = {1{$random}};
//  assign io_fpu_cp_req_bits_div = {1{$random}};
//  assign io_fpu_cp_req_bits_fma = {1{$random}};
//  assign io_fpu_cp_req_bits_fastpipe = {1{$random}};
//  assign io_fpu_cp_req_bits_toint = {1{$random}};
//  assign io_fpu_cp_req_bits_fromint = {1{$random}};
//  assign io_fpu_cp_req_bits_single = {1{$random}};
//  assign io_fpu_cp_req_bits_swap23 = {1{$random}};
//  assign io_fpu_cp_req_bits_swap12 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren3 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren2 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren1 = {1{$random}};
//  assign io_fpu_cp_req_bits_wen = {1{$random}};
//  assign io_fpu_cp_req_bits_ldst = {1{$random}};
//  assign io_fpu_cp_req_bits_cmd = {1{$random}};
//  assign io_fpu_cp_req_valid = {1{$random}};
//  assign io_imem_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T650 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T649 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign T5 = T6 | csr_io_interrupt;
  assign T6 = ctrl_killd ^ 1'h1;
  assign ctrl_killd = T7;
  assign T7 = T8 | csr_io_interrupt;
  assign T8 = T647 | ctrl_stalld;
  assign ctrl_stalld = T9 | csr_io_csr_stall;
  assign T9 = T435 | id_do_fence;
  assign id_do_fence = T60 | T10;
  assign T10 = id_mem_busy & T11;
  assign T11 = T20 | id_csr_en;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_ctrl_csr = T12;
  assign T12 = {T18, T13};
  assign T13 = {T16, T14};
  assign T14 = T15 == 32'h1070;
  assign T15 = io_imem_resp_bits_data_0 & 32'h1078;
  assign T16 = T17 == 32'h2070;
  assign T17 = io_imem_resp_bits_data_0 & 32'h2078;
  assign T18 = T19 == 32'h70;
  assign T19 = io_imem_resp_bits_data_0 & 32'h3078;
  assign T20 = T55 | T21;
  assign T21 = id_reg_fence & T22;
  assign T22 = id_ctrl_mem | id_ctrl_rocc;
  assign id_ctrl_rocc = T23;
  assign T23 = T26 | T24;
  assign T24 = T25 == 32'h58;
  assign T25 = io_imem_resp_bits_data_0 & 32'h58;
  assign T26 = T27 == 32'h8;
  assign T27 = io_imem_resp_bits_data_0 & 32'h5c;
  assign id_ctrl_mem = T28;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h1000202f;
  assign T30 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h800202f;
  assign T33 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T34 = T37 | T35;
  assign T35 = T36 == 32'h202f;
  assign T36 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'h2003;
  assign T39 = io_imem_resp_bits_data_0 & 32'h605b;
  assign T40 = T43 | T41;
  assign T41 = T42 == 32'h3;
  assign T42 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T43 = T46 | T44;
  assign T44 = T45 == 32'h3;
  assign T45 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T46 = T47 == 32'h3;
  assign T47 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T1072 = reset ? 1'h0 : T48;
  assign T48 = id_fence_next | T49;
  assign T49 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_ctrl_fence | T50;
  assign T50 = id_ctrl_amo & id_amo_rl;
  assign id_amo_rl = io_imem_resp_bits_data_0[5'h19];
  assign id_ctrl_amo = T51;
  assign T51 = T52 == 32'h200c;
  assign T52 = io_imem_resp_bits_data_0 & 32'h204c;
  assign id_ctrl_fence = T53;
  assign T53 = T54 == 32'h4;
  assign T54 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T55 = T58 | id_ctrl_fence_i;
  assign id_ctrl_fence_i = T56;
  assign T56 = T57 == 32'h1008;
  assign T57 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T58 = id_ctrl_amo & id_amo_aq;
  assign id_amo_aq = io_imem_resp_bits_data_0[5'h1a];
  assign id_mem_busy = T59 | io_dmem_req_valid;
  assign T59 = io_dmem_ordered ^ 1'h1;
  assign T60 = id_rocc_busy & id_ctrl_fence;
  assign id_rocc_busy = T431 | T61;
  assign T61 = wb_reg_valid & wb_ctrl_rocc;
  assign T62 = T650 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign T63 = T649 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign T64 = T65 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign T65 = ctrl_killd ^ 1'h1;
  assign T66 = ctrl_killm ^ 1'h1;
  assign ctrl_killm = T427 | fpu_kill_mem;
  assign fpu_kill_mem = T67 & io_fpu_nack_mem;
  assign T67 = mem_reg_valid & mem_ctrl_fp;
  assign T68 = T649 ? ex_ctrl_fp : mem_ctrl_fp;
  assign T69 = T65 ? id_ctrl_fp : ex_ctrl_fp;
  assign id_ctrl_fp = T70;
  assign T70 = T73 | T71;
  assign T71 = T72 == 32'h40;
  assign T72 = io_imem_resp_bits_data_0 & 32'h68;
  assign T73 = T76 | T74;
  assign T74 = T75 == 32'h40;
  assign T75 = io_imem_resp_bits_data_0 & 32'h70;
  assign T76 = T77 == 32'h4;
  assign T77 = io_imem_resp_bits_data_0 & 32'h5c;
  assign T78 = ctrl_killx ^ 1'h1;
  assign ctrl_killx = T81 | T79;
  assign T79 = ex_reg_valid ^ 1'h1;
  assign T80 = ctrl_killd ^ 1'h1;
  assign T81 = take_pc | replay_ex;
  assign replay_ex = ex_reg_valid & T82;
  assign T82 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T83 = T65 ? id_load_use : ex_reg_load_use;
  assign id_load_use = T84;
  assign T84 = T87 & mem_ctrl_mem;
  assign T85 = T649 ? ex_ctrl_mem : mem_ctrl_mem;
  assign T86 = T65 ? id_ctrl_mem : ex_ctrl_mem;
  assign T87 = mem_reg_valid & data_hazard_mem;
  assign data_hazard_mem = mem_ctrl_wxd & T88;
  assign T88 = T120 | T89;
  assign T89 = T91 & T90;
  assign T90 = id_waddr == mem_waddr;
  assign mem_waddr = mem_reg_inst[4'hb:3'h7];
  assign id_waddr = io_imem_resp_bits_data_0[4'hb:3'h7];
  assign T91 = id_ctrl_wxd & T92;
  assign T92 = id_waddr != 5'h0;
  assign id_ctrl_wxd = T93;
  assign T93 = T96 | T94;
  assign T94 = T95 == 32'h80000010;
  assign T95 = io_imem_resp_bits_data_0 & 32'h90000018;
  assign T96 = T99 | T97;
  assign T97 = T98 == 32'h4018;
  assign T98 = io_imem_resp_bits_data_0 & 32'h4018;
  assign T99 = T102 | T100;
  assign T100 = T101 == 32'h4000;
  assign T101 = io_imem_resp_bits_data_0 & 32'h4040;
  assign T102 = T105 | T103;
  assign T103 = T104 == 32'h2030;
  assign T104 = io_imem_resp_bits_data_0 & 32'h2038;
  assign T105 = T106 | T51;
  assign T106 = T109 | T107;
  assign T107 = T108 == 32'h1030;
  assign T108 = io_imem_resp_bits_data_0 & 32'h1038;
  assign T109 = T112 | T110;
  assign T110 = T111 == 32'h68;
  assign T111 = io_imem_resp_bits_data_0 & 32'h78;
  assign T112 = T115 | T113;
  assign T113 = T114 == 32'h24;
  assign T114 = io_imem_resp_bits_data_0 & 32'h2024;
  assign T115 = T118 | T116;
  assign T116 = T117 == 32'h10;
  assign T117 = io_imem_resp_bits_data_0 & 32'h50;
  assign T118 = T119 == 32'h0;
  assign T119 = io_imem_resp_bits_data_0 & 32'h6c;
  assign T120 = T137 | T121;
  assign T121 = T123 & T122;
  assign T122 = id_raddr_1 == mem_waddr;
  assign id_raddr_1 = io_imem_resp_bits_data_0[5'h18:5'h14];
  assign T123 = id_ctrl_rxs2 & T124;
  assign T124 = id_raddr_1 != 5'h0;
  assign id_ctrl_rxs2 = T125;
  assign T125 = T128 | T126;
  assign T126 = T127 == 32'h3018;
  assign T127 = io_imem_resp_bits_data_0 & 32'h3018;
  assign T128 = T129 | T51;
  assign T129 = T132 | T130;
  assign T130 = T131 == 32'h1008;
  assign T131 = io_imem_resp_bits_data_0 & 32'h105c;
  assign T132 = T135 | T133;
  assign T133 = T134 == 32'h30;
  assign T134 = io_imem_resp_bits_data_0 & 32'h74;
  assign T135 = T136 == 32'h20;
  assign T136 = io_imem_resp_bits_data_0 & 32'h3c;
  assign T137 = T139 & T138;
  assign T138 = id_raddr_0 == mem_waddr;
  assign id_raddr_0 = io_imem_resp_bits_data_0[5'h13:4'hf];
  assign T139 = id_ctrl_rxs1 & T140;
  assign T140 = id_raddr_0 != 5'h0;
  assign id_ctrl_rxs1 = T141;
  assign T141 = T144 | T142;
  assign T142 = T143 == 32'h0;
  assign T143 = io_imem_resp_bits_data_0 & 32'h58;
  assign T144 = T147 | T145;
  assign T145 = T146 == 32'h90000010;
  assign T146 = io_imem_resp_bits_data_0 & 32'h9000003c;
  assign T147 = T150 | T148;
  assign T148 = T149 == 32'h2018;
  assign T149 = io_imem_resp_bits_data_0 & 32'h2018;
  assign T150 = T153 | T151;
  assign T151 = T152 == 32'h2000;
  assign T152 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T153 = T156 | T154;
  assign T154 = T155 == 32'h20;
  assign T155 = io_imem_resp_bits_data_0 & 32'h38;
  assign T156 = T159 | T157;
  assign T157 = T158 == 32'h20;
  assign T158 = io_imem_resp_bits_data_0 & 32'h402c;
  assign T159 = T160 == 32'h10;
  assign T160 = io_imem_resp_bits_data_0 & 32'h54;
  assign T161 = T649 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign T162 = T65 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign wb_dcache_miss = wb_ctrl_mem & T163;
  assign T163 = io_dmem_resp_valid ^ 1'h1;
  assign T164 = T650 ? mem_ctrl_mem : wb_ctrl_mem;
  assign replay_ex_structural = T170 | T165;
  assign T165 = ex_ctrl_div & T166;
  assign T166 = div_io_req_ready ^ 1'h1;
  assign T167 = T65 ? id_ctrl_div : ex_ctrl_div;
  assign id_ctrl_div = T168;
  assign T168 = T169 == 32'h2000030;
  assign T169 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T170 = ex_ctrl_mem & T171;
  assign T171 = io_dmem_req_ready ^ 1'h1;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = T172;
  assign T172 = want_take_pc_mem & T173;
  assign T173 = mem_npc_misaligned ^ 1'h1;
  assign mem_npc_misaligned = mem_npc[1'h1];
  assign mem_npc = T174;
  assign T174 = T175 & 40'hfffffffffe;
  assign T175 = mem_ctrl_jalr ? T217 : mem_br_target;
  assign mem_br_target = T214 + T1073;
  assign T1073 = {T1077, T176};
  assign T176 = T208 ? T1074 : T177;
  assign T177 = mem_ctrl_jal ? T178 : 22'h4;
  assign T178 = T179;
  assign T179 = {T187, T180};
  assign T180 = {T183, T181};
  assign T181 = {T182, 1'h0};
  assign T182 = mem_reg_inst[5'h18:5'h15];
  assign T183 = {T185, T184};
  assign T184 = mem_reg_inst[5'h1e:5'h19];
  assign T185 = T186;
  assign T186 = mem_reg_inst[5'h14];
  assign T187 = {T191, T188};
  assign T188 = {T191, T189};
  assign T189 = T190;
  assign T190 = mem_reg_inst[5'h13:4'hc];
  assign T191 = T192;
  assign T192 = mem_reg_inst[5'h1f];
  assign T193 = T649 ? ex_ctrl_jal : mem_ctrl_jal;
  assign T194 = T65 ? id_ctrl_jal : ex_ctrl_jal;
  assign id_ctrl_jal = T110;
  assign T1074 = {T1075, T195};
  assign T195 = T196;
  assign T196 = {T204, T197};
  assign T197 = {T200, T198};
  assign T198 = {T199, 1'h0};
  assign T199 = mem_reg_inst[4'hb:4'h8];
  assign T200 = {T202, T201};
  assign T201 = mem_reg_inst[5'h1e:5'h19];
  assign T202 = T203;
  assign T203 = mem_reg_inst[3'h7];
  assign T204 = {T206, T205};
  assign T205 = {T206, T206};
  assign T206 = T207;
  assign T207 = mem_reg_inst[5'h1f];
  assign T1075 = T1076 ? 7'h7f : 7'h0;
  assign T1076 = T195[4'he];
  assign T208 = mem_ctrl_branch & mem_br_taken;
  assign mem_br_taken = bypass_mux_1[1'h0];
  assign T209 = T649 ? alu_io_out : bypass_mux_1;
  assign T210 = T649 ? ex_ctrl_branch : mem_ctrl_branch;
  assign T211 = T65 ? id_ctrl_branch : ex_ctrl_branch;
  assign id_ctrl_branch = T212;
  assign T212 = T213 == 32'h60;
  assign T213 = io_imem_resp_bits_data_0 & 32'h74;
  assign T1077 = T1078 ? 18'h3ffff : 18'h0;
  assign T1078 = T176[5'h15];
  assign T214 = mem_reg_pc;
  assign T215 = T649 ? ex_reg_pc : mem_reg_pc;
  assign T216 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T217 = T218;
  assign T218 = {T220, T219};
  assign T219 = bypass_mux_1[6'h26:1'h0];
  assign T220 = T233 ? T232 : T221;
  assign T221 = T226 ? T224 : T222;
  assign T222 = T223[1'h0];
  assign T223 = bypass_mux_1[6'h27:6'h26];
  assign T224 = T225 == 2'h3;
  assign T225 = T223;
  assign T226 = T230 | T227;
  assign T227 = T228 == 26'h3fffffe;
  assign T228 = T229;
  assign T229 = bypass_mux_1 >> 6'h26;
  assign T230 = T231 == 26'h3ffffff;
  assign T231 = T229;
  assign T232 = T223 != 2'h0;
  assign T233 = T235 | T234;
  assign T234 = T229 == 26'h1;
  assign T235 = T229 == 26'h0;
  assign T236 = T649 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign T237 = T65 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign id_ctrl_jalr = T238;
  assign T238 = T239 == 32'h24;
  assign T239 = io_imem_resp_bits_data_0 & 32'h203c;
  assign want_take_pc_mem = mem_reg_valid & T240;
  assign T240 = mem_misprediction | mem_reg_flush_pipe;
  assign T241 = T649 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign T242 = T65 ? T243 : ex_reg_flush_pipe;
  assign T243 = id_ctrl_fence_i | id_csr_flush;
  assign id_csr_flush = id_system_insn | T244;
  assign T244 = T249 & T245;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247;
  assign T247 = T248 == 12'h40;
  assign T248 = id_csr_addr & 12'h8c4;
  assign id_csr_addr = io_imem_resp_bits_data_0[5'h1f:5'h14];
  assign T249 = id_csr_en & T250;
  assign T250 = id_csr_ren ^ 1'h1;
  assign id_csr_ren = T252 & T251;
  assign T251 = id_raddr_0 == 5'h0;
  assign T252 = T254 | T253;
  assign T253 = id_ctrl_csr == 3'h3;
  assign T254 = id_ctrl_csr == 3'h2;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign mem_misprediction = T257 & T255;
  assign T255 = T256 | mem_ctrl_jal;
  assign T256 = mem_ctrl_branch | mem_ctrl_jalr;
  assign T257 = mem_wrong_npc & mem_reg_valid;
  assign mem_wrong_npc = T259 | T258;
  assign T258 = ex_reg_valid ^ 1'h1;
  assign T259 = mem_npc != ex_reg_pc;
  assign take_pc_wb = T260;
  assign T260 = T261 | csr_io_eret;
  assign T261 = replay_wb | wb_xcpt;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T262 = mem_xcpt & T263;
  assign T263 = take_pc_wb ^ 1'h1;
  assign mem_xcpt = T266 | T264;
  assign T264 = T265 & io_dmem_xcpt_pf_ld;
  assign T265 = mem_reg_valid & mem_ctrl_mem;
  assign T266 = T269 | T267;
  assign T267 = T268 & io_dmem_xcpt_pf_st;
  assign T268 = mem_reg_valid & mem_ctrl_mem;
  assign T269 = T272 | T270;
  assign T270 = T271 & io_dmem_xcpt_ma_ld;
  assign T271 = mem_reg_valid & mem_ctrl_mem;
  assign T272 = T275 | T273;
  assign T273 = T274 & io_dmem_xcpt_ma_st;
  assign T274 = mem_reg_valid & mem_ctrl_mem;
  assign T275 = T277 | T276;
  assign T276 = want_take_pc_mem & mem_npc_misaligned;
  assign T277 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T278 = T415 & ex_xcpt;
  assign ex_xcpt = T280 | T279;
  assign T279 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign T280 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T281 = T411 & id_xcpt;
  assign id_xcpt = T410 | id_illegal_insn;
  assign id_illegal_insn = T285 | T282;
  assign T282 = id_ctrl_rocc & T283;
  assign T283 = T284 ^ 1'h1;
  assign T284 = csr_io_status_xs != 2'h0;
  assign T285 = T289 | T286;
  assign T286 = id_ctrl_fp & T287;
  assign T287 = T288 ^ 1'h1;
  assign T288 = csr_io_status_fs != 2'h0;
  assign T289 = id_ctrl_legal ^ 1'h1;
  assign id_ctrl_legal = T290;
  assign T290 = T293 | T291;
  assign T291 = T292 == 32'h3;
  assign T292 = io_imem_resp_bits_data_0 & 32'h7067;
  assign T293 = T296 | T294;
  assign T294 = T295 == 32'h33;
  assign T295 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T296 = T299 | T297;
  assign T297 = T298 == 32'h4063;
  assign T298 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T299 = T302 | T300;
  assign T300 = T301 == 32'h1063;
  assign T301 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T302 = T305 | T303;
  assign T303 = T304 == 32'h23;
  assign T304 = io_imem_resp_bits_data_0 & 32'h603f;
  assign T305 = T308 | T306;
  assign T306 = T307 == 32'he0000053;
  assign T307 = io_imem_resp_bits_data_0 & 32'hedf0707f;
  assign T308 = T311 | T309;
  assign T309 = T310 == 32'he0000053;
  assign T310 = io_imem_resp_bits_data_0 & 32'hfdf0607f;
  assign T311 = T314 | T312;
  assign T312 = T313 == 32'hc0000053;
  assign T313 = io_imem_resp_bits_data_0 & 32'hedc0007f;
  assign T314 = T317 | T315;
  assign T315 = T316 == 32'h58000053;
  assign T316 = io_imem_resp_bits_data_0 & 32'hfdf0007f;
  assign T317 = T320 | T318;
  assign T318 = T319 == 32'h42000053;
  assign T319 = io_imem_resp_bits_data_0 & 32'h7ff0007f;
  assign T320 = T323 | T321;
  assign T321 = T322 == 32'h40100053;
  assign T322 = io_imem_resp_bits_data_0 & 32'h7ff0007f;
  assign T323 = T325 | T324;
  assign T324 = io_imem_resp_bits_data_0 == 32'h30500073;
  assign T325 = T328 | T326;
  assign T326 = T327 == 32'h20000053;
  assign T327 = io_imem_resp_bits_data_0 & 32'h7c00507f;
  assign T328 = T331 | T329;
  assign T329 = T330 == 32'h20000053;
  assign T330 = io_imem_resp_bits_data_0 & 32'h7c00607f;
  assign T331 = T334 | T332;
  assign T332 = T333 == 32'h20000053;
  assign T333 = io_imem_resp_bits_data_0 & 32'hf400607f;
  assign T334 = T337 | T335;
  assign T335 = T336 == 32'h10100073;
  assign T336 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T337 = T338 | T29;
  assign T338 = T341 | T339;
  assign T339 = T340 == 32'h10000073;
  assign T340 = io_imem_resp_bits_data_0 & 32'hffdfffff;
  assign T341 = T342 | T32;
  assign T342 = T345 | T343;
  assign T343 = T344 == 32'h2004033;
  assign T344 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T345 = T348 | T346;
  assign T346 = T347 == 32'h5033;
  assign T347 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T348 = T351 | T349;
  assign T349 = T350 == 32'h501b;
  assign T350 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T351 = T354 | T352;
  assign T352 = T353 == 32'h5013;
  assign T353 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T354 = T357 | T355;
  assign T355 = T356 == 32'h2073;
  assign T356 = io_imem_resp_bits_data_0 & 32'h2077;
  assign T357 = T360 | T358;
  assign T358 = T359 == 32'h205b;
  assign T359 = io_imem_resp_bits_data_0 & 32'h205f;
  assign T360 = T361 | T35;
  assign T361 = T364 | T362;
  assign T362 = T363 == 32'h2013;
  assign T363 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T364 = T367 | T365;
  assign T365 = T366 == 32'h200b;
  assign T366 = io_imem_resp_bits_data_0 & 32'h205f;
  assign T367 = T368 | T38;
  assign T368 = T371 | T369;
  assign T369 = T370 == 32'h101b;
  assign T370 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T371 = T374 | T372;
  assign T372 = T373 == 32'h1013;
  assign T373 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T374 = T377 | T375;
  assign T375 = T376 == 32'h73;
  assign T376 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T377 = T380 | T378;
  assign T378 = T379 == 32'h6f;
  assign T379 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T380 = T383 | T381;
  assign T381 = T382 == 32'h63;
  assign T382 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T383 = T386 | T384;
  assign T384 = T385 == 32'h5b;
  assign T385 = io_imem_resp_bits_data_0 & 32'h105f;
  assign T386 = T389 | T387;
  assign T387 = T388 == 32'h53;
  assign T388 = io_imem_resp_bits_data_0 & 32'he400007f;
  assign T389 = T392 | T390;
  assign T390 = T391 == 32'h43;
  assign T391 = io_imem_resp_bits_data_0 & 32'h4000073;
  assign T392 = T395 | T393;
  assign T393 = T394 == 32'h33;
  assign T394 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T395 = T398 | T396;
  assign T396 = T397 == 32'h33;
  assign T397 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T398 = T401 | T399;
  assign T399 = T400 == 32'h17;
  assign T400 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T401 = T404 | T402;
  assign T402 = T403 == 32'hf;
  assign T403 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T404 = T407 | T405;
  assign T405 = T406 == 32'hb;
  assign T406 = io_imem_resp_bits_data_0 & 32'h105f;
  assign T407 = T44 | T408;
  assign T408 = T409 == 32'h3;
  assign T409 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T410 = csr_io_interrupt | io_imem_resp_bits_xcpt_if;
  assign T411 = ctrl_killd ^ 1'h1;
  assign T412 = T413 & io_imem_resp_valid;
  assign T413 = csr_io_interrupt & T414;
  assign T414 = take_pc ^ 1'h1;
  assign T415 = ctrl_killx ^ 1'h1;
  assign T416 = T417 & ex_reg_xcpt_interrupt;
  assign T417 = take_pc ^ 1'h1;
  assign replay_wb = replay_wb_common | T418;
  assign T418 = T420 & T419;
  assign T419 = io_rocc_cmd_ready ^ 1'h1;
  assign T420 = wb_reg_valid & wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T421 = replay_mem & T422;
  assign T422 = take_pc_wb ^ 1'h1;
  assign replay_mem = T423 | fpu_kill_mem;
  assign T423 = dcache_kill_mem | mem_reg_replay;
  assign T424 = T425 & replay_ex;
  assign T425 = take_pc ^ 1'h1;
  assign dcache_kill_mem = T426 & io_dmem_replay_next_valid;
  assign T426 = mem_reg_valid & mem_ctrl_wxd;
  assign T427 = killm_common | mem_xcpt;
  assign killm_common = T429 | T428;
  assign T428 = mem_reg_valid ^ 1'h1;
  assign T429 = T430 | mem_reg_xcpt;
  assign T430 = dcache_kill_mem | take_pc_wb;
  assign T431 = T433 | T432;
  assign T432 = mem_reg_valid & mem_ctrl_rocc;
  assign T433 = io_rocc_busy | T434;
  assign T434 = ex_reg_valid & ex_ctrl_rocc;
  assign T435 = T444 | T436;
  assign T436 = T438 & T437;
  assign T437 = io_rocc_cmd_ready ^ 1'h1;
  assign T438 = wb_reg_rocc_pending & id_ctrl_rocc;
  assign T1079 = reset ? 1'h0 : T439;
  assign T439 = wb_reg_xcpt ? 1'h0 : T440;
  assign T440 = wb_rocc_val ? T441 : wb_reg_rocc_pending;
  assign T441 = io_rocc_cmd_ready ^ 1'h1;
  assign wb_rocc_val = T443 & T442;
  assign T442 = replay_wb_common ^ 1'h1;
  assign T443 = wb_reg_valid & wb_ctrl_rocc;
  assign T444 = T447 | T445;
  assign T445 = id_ctrl_mem & T446;
  assign T446 = io_dmem_req_ready ^ 1'h1;
  assign T447 = T500 | T448;
  assign T448 = id_ctrl_fp & id_stall_fpu;
  assign id_stall_fpu = T498 | T449;
  assign T449 = T490 | T450;
  assign T450 = io_fpu_dec_wen & T451;
  assign T451 = R452[id_waddr];
  assign T1080 = reset ? 32'h0 : T453;
  assign T453 = T489 ? T485 : T454;
  assign T454 = T484 ? T477 : T455;
  assign T455 = T459 ? T456 : R452;
  assign T456 = R452 | T457;
  assign T457 = T459 ? T458 : 32'h0;
  assign T458 = 1'h1 << wb_waddr;
  assign wb_waddr = wb_reg_inst[4'hb:3'h7];
  assign T459 = T463 & wb_valid;
  assign wb_valid = T461 & T460;
  assign T460 = csr_io_csr_xcpt ^ 1'h1;
  assign T461 = wb_reg_valid & T462;
  assign T462 = replay_wb ^ 1'h1;
  assign T463 = T464 | io_fpu_sboard_set;
  assign T464 = wb_dcache_miss & wb_ctrl_wfd;
  assign T465 = T650 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign T466 = T649 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign T467 = T65 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign id_ctrl_wfd = T468;
  assign T468 = T471 | T469;
  assign T469 = T470 == 32'h10000040;
  assign T470 = io_imem_resp_bits_data_0 & 32'h10000068;
  assign T471 = T472 | T74;
  assign T472 = T475 | T473;
  assign T473 = T474 == 32'h40;
  assign T474 = io_imem_resp_bits_data_0 & 32'h80000068;
  assign T475 = T476 == 32'h4;
  assign T476 = io_imem_resp_bits_data_0 & 32'h3c;
  assign T477 = T456 & T478;
  assign T478 = ~ T479;
  assign T479 = T482 ? T480 : 32'h0;
  assign T480 = 1'h1 << dmem_resp_waddr;
  assign dmem_resp_waddr = T481[3'h5:1'h1];
  assign T481 = io_dmem_resp_bits_tag;
  assign T482 = dmem_resp_replay & dmem_resp_fpu;
  assign dmem_resp_fpu = T483;
  assign T483 = io_dmem_resp_bits_tag[1'h0];
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T484 = T459 | T482;
  assign T485 = T477 & T486;
  assign T486 = ~ T487;
  assign T487 = io_fpu_sboard_clr ? T488 : 32'h0;
  assign T488 = 1'h1 << io_fpu_sboard_clra;
  assign T489 = T484 | io_fpu_sboard_clr;
  assign T490 = T493 | T491;
  assign T491 = io_fpu_dec_ren3 & T492;
  assign T492 = R452[id_raddr3];
  assign id_raddr3 = io_imem_resp_bits_data_0[5'h1f:5'h1b];
  assign T493 = T496 | T494;
  assign T494 = io_fpu_dec_ren2 & T495;
  assign T495 = R452[id_raddr_1];
  assign T496 = io_fpu_dec_ren1 & T497;
  assign T497 = R452[id_raddr_0];
  assign T498 = id_csr_en & T499;
  assign T499 = io_fpu_fcsr_rdy ^ 1'h1;
  assign T500 = T533 | id_sboard_hazard;
  assign id_sboard_hazard = T528 | T501;
  assign T501 = T91 & T502;
  assign T502 = T503[id_waddr];
  assign T503 = R516 & T504;
  assign T504 = ~ T505;
  assign T505 = ll_wen ? T506 : 32'h0;
  assign T506 = 1'h1 << ll_waddr;
  assign ll_waddr = T507;
  assign T507 = T510 ? dmem_resp_waddr : T508;
  assign T508 = T509 ? io_rocc_resp_bits_rd : div_io_resp_bits_tag;
  assign T509 = io_rocc_resp_ready & io_rocc_resp_valid;
  assign T510 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_xpu = T511 ^ 1'h1;
  assign T511 = T512;
  assign T512 = io_dmem_resp_bits_tag[1'h0];
  assign ll_wen = T513;
  assign T513 = T510 ? 1'h1 : T514;
  assign T514 = T509 ? 1'h1 : T515;
  assign T515 = T770 & div_io_resp_valid;
  assign T1081 = reset ? 32'h0 : T517;
  assign T517 = T527 ? T519 : T518;
  assign T518 = ll_wen ? T503 : R516;
  assign T519 = T503 | T520;
  assign T520 = T522 ? T521 : 32'h0;
  assign T521 = 1'h1 << wb_waddr;
  assign T522 = wb_set_sboard & wb_wen;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign T523 = T650 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign wb_set_sboard = T524 | wb_ctrl_rocc;
  assign T524 = wb_ctrl_div | wb_dcache_miss;
  assign T525 = T650 ? mem_ctrl_div : wb_ctrl_div;
  assign T526 = T649 ? ex_ctrl_div : mem_ctrl_div;
  assign T527 = ll_wen | T522;
  assign T528 = T531 | T529;
  assign T529 = T123 & T530;
  assign T530 = T503[id_raddr_1];
  assign T531 = T139 & T532;
  assign T532 = T503[id_raddr_0];
  assign T533 = T555 | id_wb_hazard;
  assign id_wb_hazard = wb_reg_valid & T534;
  assign T534 = T546 | fp_data_hazard_wb;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T535;
  assign T535 = T538 | T536;
  assign T536 = io_fpu_dec_wen & T537;
  assign T537 = id_waddr == wb_waddr;
  assign T538 = T541 | T539;
  assign T539 = io_fpu_dec_ren3 & T540;
  assign T540 = id_raddr3 == wb_waddr;
  assign T541 = T544 | T542;
  assign T542 = io_fpu_dec_ren2 & T543;
  assign T543 = id_raddr_1 == wb_waddr;
  assign T544 = io_fpu_dec_ren1 & T545;
  assign T545 = id_raddr_0 == wb_waddr;
  assign T546 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_ctrl_wxd & T547;
  assign T547 = T550 | T548;
  assign T548 = T91 & T549;
  assign T549 = id_waddr == wb_waddr;
  assign T550 = T553 | T551;
  assign T551 = T123 & T552;
  assign T552 = id_raddr_1 == wb_waddr;
  assign T553 = T139 & T554;
  assign T554 = id_raddr_0 == wb_waddr;
  assign T555 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = mem_reg_valid & T556;
  assign T556 = T568 | fp_data_hazard_mem;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T557;
  assign T557 = T560 | T558;
  assign T558 = io_fpu_dec_wen & T559;
  assign T559 = id_waddr == mem_waddr;
  assign T560 = T563 | T561;
  assign T561 = io_fpu_dec_ren3 & T562;
  assign T562 = id_raddr3 == mem_waddr;
  assign T563 = T566 | T564;
  assign T564 = io_fpu_dec_ren2 & T565;
  assign T565 = id_raddr_1 == mem_waddr;
  assign T566 = io_fpu_dec_ren1 & T567;
  assign T567 = id_raddr_0 == mem_waddr;
  assign T568 = data_hazard_mem & mem_cannot_bypass;
  assign mem_cannot_bypass = T569 | mem_ctrl_rocc;
  assign T569 = T570 | mem_ctrl_fp;
  assign T570 = T571 | mem_ctrl_div;
  assign T571 = T617 | T572;
  assign T572 = mem_ctrl_mem & mem_mem_cmd_bh;
  assign T573 = T649 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T590 | T574;
  assign T574 = T585 | T575;
  assign T575 = 3'h5 == ex_ctrl_mem_type;
  assign T576 = T65 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign id_ctrl_mem_type = T577;
  assign T577 = {T583, T578};
  assign T578 = {T581, T579};
  assign T579 = T580 == 32'h1000;
  assign T580 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T581 = T582 == 32'h2000;
  assign T582 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T583 = T584 == 32'h4000;
  assign T584 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T585 = T587 | T586;
  assign T586 = 3'h1 == ex_ctrl_mem_type;
  assign T587 = T589 | T588;
  assign T588 = 3'h4 == ex_ctrl_mem_type;
  assign T589 = 3'h0 == ex_ctrl_mem_type;
  assign T590 = ex_ctrl_mem_cmd == 5'h7;
  assign T591 = T65 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign id_ctrl_mem_cmd = T592;
  assign T592 = {1'h0, T593};
  assign T593 = {T615, T594};
  assign T594 = {T609, T595};
  assign T595 = {T604, T596};
  assign T596 = T599 | T597;
  assign T597 = T598 == 32'h20000020;
  assign T598 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T599 = T602 | T600;
  assign T600 = T601 == 32'h18000020;
  assign T601 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T602 = T603 == 32'h20;
  assign T603 = io_imem_resp_bits_data_0 & 32'h28;
  assign T604 = T607 | T605;
  assign T605 = T606 == 32'h40000008;
  assign T606 = io_imem_resp_bits_data_0 & 32'h40000008;
  assign T607 = T608 == 32'h10000008;
  assign T608 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T609 = T612 | T610;
  assign T610 = T611 == 32'h80000008;
  assign T611 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T612 = T613 | T607;
  assign T613 = T614 == 32'h8000008;
  assign T614 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T615 = T616 == 32'h8;
  assign T616 = io_imem_resp_bits_data_0 & 32'h18000008;
  assign T617 = mem_ctrl_csr != 3'h0;
  assign T618 = T649 ? ex_ctrl_csr : mem_ctrl_csr;
  assign T619 = T65 ? id_csr : T620;
  assign T620 = T65 ? id_ctrl_csr : ex_ctrl_csr;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_ex_hazard = ex_reg_valid & T621;
  assign T621 = T633 | fp_data_hazard_ex;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T622;
  assign T622 = T625 | T623;
  assign T623 = io_fpu_dec_wen & T624;
  assign T624 = id_waddr == ex_waddr;
  assign ex_waddr = ex_reg_inst[4'hb:3'h7];
  assign T625 = T628 | T626;
  assign T626 = io_fpu_dec_ren3 & T627;
  assign T627 = id_raddr3 == ex_waddr;
  assign T628 = T631 | T629;
  assign T629 = io_fpu_dec_ren2 & T630;
  assign T630 = id_raddr_1 == ex_waddr;
  assign T631 = io_fpu_dec_ren1 & T632;
  assign T632 = id_raddr_0 == ex_waddr;
  assign T633 = data_hazard_ex & ex_cannot_bypass;
  assign ex_cannot_bypass = T634 | ex_ctrl_rocc;
  assign T634 = T635 | ex_ctrl_fp;
  assign T635 = T636 | ex_ctrl_div;
  assign T636 = T637 | ex_ctrl_mem;
  assign T637 = T638 | ex_ctrl_jalr;
  assign T638 = ex_ctrl_csr != 3'h0;
  assign data_hazard_ex = ex_ctrl_wxd & T639;
  assign T639 = T642 | T640;
  assign T640 = T91 & T641;
  assign T641 = id_waddr == ex_waddr;
  assign T642 = T645 | T643;
  assign T643 = T123 & T644;
  assign T644 = id_raddr_1 == ex_waddr;
  assign T645 = T139 & T646;
  assign T646 = id_raddr_0 == ex_waddr;
  assign T647 = T648 | take_pc;
  assign T648 = io_imem_resp_valid ^ 1'h1;
  assign T649 = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T650 = T651 | mem_reg_xcpt_interrupt;
  assign T651 = mem_reg_valid | mem_reg_replay;
  assign T652 = wb_reg_inst;
  assign T653 = R654;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T708 : T656;
  assign T656 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T657 = T697 ? T671 : T658;
  assign T658 = T65 ? T659 : ex_reg_rs_lsb_1;
  assign T659 = T670 ? 2'h0 : T660;
  assign T660 = T667 ? 2'h1 : T661;
  assign T661 = T662 ? 2'h2 : 2'h3;
  assign T662 = T664 & T663;
  assign T663 = mem_waddr == id_raddr_1;
  assign T664 = T666 & T665;
  assign T665 = mem_ctrl_mem ^ 1'h1;
  assign T666 = mem_reg_valid & mem_ctrl_wxd;
  assign T667 = T669 & T668;
  assign T668 = ex_waddr == id_raddr_1;
  assign T669 = ex_reg_valid & ex_ctrl_wxd;
  assign T670 = 5'h0 == id_raddr_1;
  assign T671 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T672;
  assign T672 = T695 ? rf_wdata : T673;
  assign T673 = T674[T682];
  assign T676 = T679 & T677;
  assign T677 = T678 < 5'h1f;
  assign T678 = T681;
  assign T679 = rf_wen & T680;
  assign T680 = rf_waddr != 5'h0;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign rf_wen = wb_wen | ll_wen;
  assign T681 = ~ rf_waddr;
  assign T682 = ~ T683;
  assign T683 = id_raddr_1;
  assign rf_wdata = T694 ? io_dmem_resp_bits_data : T684;
  assign T684 = ll_wen ? ll_wdata : T685;
  assign T685 = T691 ? csr_io_rw_rdata : bypass_mux_2;
  assign T686 = T650 ? T687 : bypass_mux_2;
  assign T687 = T690 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = T688;
  assign T688 = mem_ctrl_jalr ? T1082 : T689;
  assign T689 = bypass_mux_1;
  assign T1082 = {T1083, mem_br_target};
  assign T1083 = T1084 ? 24'hffffff : 24'h0;
  assign T1084 = mem_br_target[6'h27];
  assign T690 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T691 = wb_ctrl_csr != 3'h0;
  assign T692 = T650 ? mem_ctrl_csr : wb_ctrl_csr;
  assign ll_wdata = T693;
  assign T693 = T509 ? io_rocc_resp_bits_data : div_io_resp_bits_data;
  assign T694 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T695 = T679 & T696;
  assign T696 = rf_waddr == id_raddr_1;
  assign T697 = T65 & T698;
  assign T698 = id_ctrl_rxs2 & T699;
  assign T699 = T700 ^ 1'h1;
  assign T700 = T704 | T701;
  assign T701 = T703 & T702;
  assign T702 = mem_waddr == id_raddr_1;
  assign T703 = mem_reg_valid & mem_ctrl_wxd;
  assign T704 = T705 | T662;
  assign T705 = T670 | T667;
  assign T706 = T697 ? T707 : ex_reg_rs_msb_1;
  assign T707 = id_rs_1 >> 2'h2;
  assign T708 = T714 ? T712 : T709;
  assign T709 = T710 ? bypass_mux_1 : 64'h0;
  assign T710 = T711[1'h0];
  assign T711 = ex_reg_rs_lsb_1;
  assign T712 = T713 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T713 = T711[1'h0];
  assign T714 = T711[1'h1];
  assign T715 = T65 ? T700 : ex_reg_rs_bypass_1;
  assign T716 = T717;
  assign T717 = wb_reg_inst[5'h18:5'h14];
  assign T718 = R719;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T749 : T721;
  assign T721 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T722 = T739 ? T732 : T723;
  assign T723 = T65 ? T724 : ex_reg_rs_lsb_0;
  assign T724 = T731 ? 2'h0 : T725;
  assign T725 = T729 ? 2'h1 : T726;
  assign T726 = T727 ? 2'h2 : 2'h3;
  assign T727 = T664 & T728;
  assign T728 = mem_waddr == id_raddr_0;
  assign T729 = T669 & T730;
  assign T730 = ex_waddr == id_raddr_0;
  assign T731 = 5'h0 == id_raddr_0;
  assign T732 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T733;
  assign T733 = T737 ? rf_wdata : T734;
  assign T734 = T674[T735];
  assign T735 = ~ T736;
  assign T736 = id_raddr_0;
  assign T737 = T679 & T738;
  assign T738 = rf_waddr == id_raddr_0;
  assign T739 = T65 & T740;
  assign T740 = id_ctrl_rxs1 & T741;
  assign T741 = T742 ^ 1'h1;
  assign T742 = T745 | T743;
  assign T743 = T703 & T744;
  assign T744 = mem_waddr == id_raddr_0;
  assign T745 = T746 | T727;
  assign T746 = T731 | T729;
  assign T747 = T739 ? T748 : ex_reg_rs_msb_0;
  assign T748 = id_rs_0 >> 2'h2;
  assign T749 = T755 ? T753 : T750;
  assign T750 = T751 ? bypass_mux_1 : 64'h0;
  assign T751 = T752[1'h0];
  assign T752 = ex_reg_rs_lsb_0;
  assign T753 = T754 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T754 = T752[1'h0];
  assign T755 = T752[1'h1];
  assign T756 = T65 ? T742 : ex_reg_rs_bypass_0;
  assign T757 = T758;
  assign T758 = wb_reg_inst[5'h13:4'hf];
  assign T759 = rf_wen;
  assign T760 = rf_wdata;
  assign T761 = T762;
  assign T762 = rf_wen ? rf_waddr : 5'h0;
  assign T763 = wb_reg_pc;
  assign T764 = T650 ? mem_reg_pc : wb_reg_pc;
  assign T765 = wb_valid;
  assign T766 = T767;
  assign T767 = csr_io_time[6'h20:1'h0];
  assign T768 = io_host_id;
  assign T770 = T510 ? 1'h0 : T771;
  assign T771 = T509 ? 1'h0 : T772;
  assign T772 = T773 ^ 1'h1;
  assign T773 = wb_reg_valid & wb_ctrl_wxd;
  assign T774 = killm_common & R775;
  assign T776 = div_io_req_ready & T833;
  assign T777 = T65 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign id_ctrl_alu_dw = T778;
  assign T778 = T781 | T779;
  assign T779 = T780 == 32'h40;
  assign T780 = io_imem_resp_bits_data_0 & 32'h40;
  assign T781 = T784 | T782;
  assign T782 = T783 == 32'h0;
  assign T783 = io_imem_resp_bits_data_0 & 32'h8;
  assign T784 = T785 == 32'h0;
  assign T785 = io_imem_resp_bits_data_0 & 32'h10;
  assign T786 = T65 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign id_ctrl_alu_fn = T787;
  assign T787 = {T826, T788};
  assign T788 = {T815, T789};
  assign T789 = {T798, T790};
  assign T790 = T793 | T791;
  assign T791 = T792 == 32'h5010;
  assign T792 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T793 = T796 | T794;
  assign T794 = T795 == 32'h1040;
  assign T795 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T796 = T797 == 32'h1010;
  assign T797 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T798 = T801 | T799;
  assign T799 = T800 == 32'h40001010;
  assign T800 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T801 = T804 | T802;
  assign T802 = T803 == 32'h40000030;
  assign T803 = io_imem_resp_bits_data_0 & 32'h40000074;
  assign T804 = T807 | T805;
  assign T805 = T806 == 32'h6010;
  assign T806 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T807 = T810 | T808;
  assign T808 = T809 == 32'h3010;
  assign T809 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T810 = T813 | T811;
  assign T811 = T812 == 32'h2040;
  assign T812 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T813 = T814 == 32'h40;
  assign T814 = io_imem_resp_bits_data_0 & 32'h4054;
  assign T815 = T818 | T816;
  assign T816 = T817 == 32'h4040;
  assign T817 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T818 = T821 | T819;
  assign T819 = T820 == 32'h4010;
  assign T820 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T821 = T824 | T822;
  assign T822 = T823 == 32'h4010;
  assign T823 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T824 = T825 == 32'h2010;
  assign T825 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T826 = T829 | T827;
  assign T827 = T828 == 32'h40001010;
  assign T828 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T829 = T830 | T802;
  assign T830 = T831 | T816;
  assign T831 = T832 == 32'h2010;
  assign T832 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T833 = ex_reg_valid & ex_ctrl_div;
  assign T834 = ex_op1;
  assign ex_op1 = T863 ? T862 : T1085;
  assign T1085 = {T1086, T835};
  assign T835 = T837 ? T836 : 40'h0;
  assign T836 = ex_reg_pc;
  assign T837 = ex_ctrl_sel_alu1 == 2'h2;
  assign T838 = T65 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign id_ctrl_sel_alu1 = T839;
  assign T839 = {T857, T840};
  assign T840 = T843 | T841;
  assign T841 = T842 == 32'h8;
  assign T842 = io_imem_resp_bits_data_0 & 32'hc;
  assign T843 = T846 | T844;
  assign T844 = T845 == 32'h0;
  assign T845 = io_imem_resp_bits_data_0 & 32'h18;
  assign T846 = T849 | T847;
  assign T847 = T848 == 32'h0;
  assign T848 = io_imem_resp_bits_data_0 & 32'h24;
  assign T849 = T852 | T850;
  assign T850 = T851 == 32'h0;
  assign T851 = io_imem_resp_bits_data_0 & 32'h44;
  assign T852 = T855 | T853;
  assign T853 = T854 == 32'h0;
  assign T854 = io_imem_resp_bits_data_0 & 32'h50;
  assign T855 = T856 == 32'h0;
  assign T856 = io_imem_resp_bits_data_0 & 32'h4004;
  assign T857 = T860 | T858;
  assign T858 = T859 == 32'h48;
  assign T859 = io_imem_resp_bits_data_0 & 32'h58;
  assign T860 = T861 == 32'h14;
  assign T861 = io_imem_resp_bits_data_0 & 32'h34;
  assign T1086 = T1087 ? 24'hffffff : 24'h0;
  assign T1087 = T835[6'h27];
  assign T862 = ex_rs_0;
  assign T863 = ex_ctrl_sel_alu1 == 2'h1;
  assign T864 = ex_op2;
  assign ex_op2 = T962 ? T961 : T1088;
  assign T1088 = {T1094, T865};
  assign T865 = T960 ? ex_imm : T1089;
  assign T1089 = {T1090, T866};
  assign T866 = T867 ? 4'h4 : 4'h0;
  assign T867 = ex_ctrl_sel_alu2 == 2'h1;
  assign T868 = T65 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign id_ctrl_sel_alu2 = T869;
  assign T869 = {T880, T870};
  assign T870 = T873 | T871;
  assign T871 = T872 == 32'h4050;
  assign T872 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T873 = T874 | T858;
  assign T874 = T877 | T875;
  assign T875 = T876 == 32'h10;
  assign T876 = io_imem_resp_bits_data_0 & 32'h70;
  assign T877 = T142 | T878;
  assign T878 = T879 == 32'h4;
  assign T879 = io_imem_resp_bits_data_0 & 32'hc;
  assign T880 = T883 | T881;
  assign T881 = T882 == 32'h4000;
  assign T882 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T883 = T844 | T116;
  assign T1090 = T1091 ? 28'hfffffff : 28'h0;
  assign T1091 = T866[2'h3];
  assign ex_imm = T884;
  assign T884 = {T948, T885};
  assign T885 = {T926, T886};
  assign T886 = {T915, T887};
  assign T887 = T914 ? T913 : T888;
  assign T888 = T912 ? T911 : T889;
  assign T889 = T891 ? T890 : 1'h0;
  assign T890 = ex_reg_inst[4'hf];
  assign T891 = ex_ctrl_sel_imm == 3'h5;
  assign T892 = T65 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign id_ctrl_sel_imm = T893;
  assign T893 = {T903, T894};
  assign T894 = {T900, T895};
  assign T895 = T898 | T896;
  assign T896 = T897 == 32'h40;
  assign T897 = io_imem_resp_bits_data_0 & 32'h44;
  assign T898 = T899 == 32'h8;
  assign T899 = io_imem_resp_bits_data_0 & 32'h18;
  assign T900 = T898 | T901;
  assign T901 = T902 == 32'h14;
  assign T902 = io_imem_resp_bits_data_0 & 32'h14;
  assign T903 = T906 | T904;
  assign T904 = T905 == 32'h10;
  assign T905 = io_imem_resp_bits_data_0 & 32'h14;
  assign T906 = T909 | T907;
  assign T907 = T908 == 32'h4;
  assign T908 = io_imem_resp_bits_data_0 & 32'h201c;
  assign T909 = T910 == 32'h0;
  assign T910 = io_imem_resp_bits_data_0 & 32'h30;
  assign T911 = ex_reg_inst[5'h14];
  assign T912 = ex_ctrl_sel_imm == 3'h4;
  assign T913 = ex_reg_inst[3'h7];
  assign T914 = ex_ctrl_sel_imm == 3'h0;
  assign T915 = T925 ? 4'h0 : T916;
  assign T916 = T922 ? T921 : T917;
  assign T917 = T920 ? T919 : T918;
  assign T918 = ex_reg_inst[5'h18:5'h15];
  assign T919 = ex_reg_inst[5'h13:5'h10];
  assign T920 = ex_ctrl_sel_imm == 3'h5;
  assign T921 = ex_reg_inst[4'hb:4'h8];
  assign T922 = T924 | T923;
  assign T923 = ex_ctrl_sel_imm == 3'h1;
  assign T924 = ex_ctrl_sel_imm == 3'h0;
  assign T925 = ex_ctrl_sel_imm == 3'h2;
  assign T926 = {T932, T927};
  assign T927 = T929 ? 6'h0 : T928;
  assign T928 = ex_reg_inst[5'h1e:5'h19];
  assign T929 = T931 | T930;
  assign T930 = ex_ctrl_sel_imm == 3'h5;
  assign T931 = ex_ctrl_sel_imm == 3'h2;
  assign T932 = T945 ? 1'h0 : T933;
  assign T933 = T944 ? T942 : T934;
  assign T934 = T941 ? T939 : T935;
  assign T935 = T938 ? 1'h0 : T936;
  assign T936 = T937;
  assign T937 = ex_reg_inst[5'h1f];
  assign T938 = ex_ctrl_sel_imm == 3'h5;
  assign T939 = T940;
  assign T940 = ex_reg_inst[3'h7];
  assign T941 = ex_ctrl_sel_imm == 3'h1;
  assign T942 = T943;
  assign T943 = ex_reg_inst[5'h14];
  assign T944 = ex_ctrl_sel_imm == 3'h3;
  assign T945 = T947 | T946;
  assign T946 = ex_ctrl_sel_imm == 3'h5;
  assign T947 = ex_ctrl_sel_imm == 3'h2;
  assign T948 = {T935, T949};
  assign T949 = {T956, T950};
  assign T950 = T953 ? T1092 : T951;
  assign T951 = T952;
  assign T952 = ex_reg_inst[5'h13:4'hc];
  assign T1092 = T935 ? 8'hff : 8'h0;
  assign T953 = T955 & T954;
  assign T954 = ex_ctrl_sel_imm != 3'h3;
  assign T955 = ex_ctrl_sel_imm != 3'h2;
  assign T956 = T959 ? T957 : T1093;
  assign T1093 = T935 ? 11'h7ff : 11'h0;
  assign T957 = T958;
  assign T958 = ex_reg_inst[5'h1e:5'h14];
  assign T959 = ex_ctrl_sel_imm == 3'h2;
  assign T960 = ex_ctrl_sel_alu2 == 2'h3;
  assign T1094 = T1095 ? 32'hffffffff : 32'h0;
  assign T1095 = T865[5'h1f];
  assign T961 = ex_rs_1;
  assign T962 = ex_ctrl_sel_alu2 == 2'h2;
  assign T963 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T277 ? mem_reg_cause : T1096;
  assign T1096 = {61'h0, T964};
  assign T964 = T276 ? 3'h0 : T965;
  assign T965 = T273 ? 3'h6 : T966;
  assign T966 = T270 ? 3'h4 : T967;
  assign T967 = T267 ? 3'h7 : 3'h5;
  assign T968 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T280 ? ex_reg_cause : 64'h2;
  assign T969 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : T1097;
  assign T1097 = {62'h0, T970};
  assign T970 = io_imem_resp_bits_xcpt_if ? 2'h1 : 2'h2;
  assign T971 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T972 = wb_reg_inst[5'h1f:5'h14];
  assign io_rocc_csr_wen = csr_io_rocc_csr_wen;
  assign io_rocc_csr_wdata = csr_io_rocc_csr_wdata;
  assign io_rocc_csr_waddr = csr_io_rocc_csr_waddr;
  assign io_rocc_exception = T973;
  assign T973 = wb_xcpt & T974;
  assign T974 = csr_io_status_xs != 2'h0;
  assign io_rocc_s = T975;
  assign T975 = csr_io_status_prv != 2'h0;
  assign io_rocc_resp_ready = T976;
  assign T976 = T510 ? 1'h0 : T977;
  assign T977 = T978 ^ 1'h1;
  assign T978 = wb_reg_valid & wb_ctrl_wxd;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T979 = T985 ? mem_reg_rs2 : wb_reg_rs2;
  assign T980 = T981 ? ex_rs_1 : mem_reg_rs2;
  assign T981 = T649 & T982;
  assign T982 = ex_ctrl_rxs2 & T983;
  assign T983 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T984 = T65 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign T985 = T650 & mem_ctrl_rocc;
  assign io_rocc_cmd_bits_rs1 = bypass_mux_2;
  assign io_rocc_cmd_bits_inst_opcode = T986;
  assign T986 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T987;
  assign T987 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T988;
  assign T988 = wb_reg_inst[4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T989;
  assign T989 = wb_reg_inst[4'hd];
  assign io_rocc_cmd_bits_inst_xd = T990;
  assign T990 = wb_reg_inst[4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T991;
  assign T991 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T992;
  assign T992 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T993;
  assign T993 = wb_reg_inst[5'h1f:5'h19];
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T994;
  assign T994 = T995 & id_ctrl_fp;
  assign T995 = ctrl_killd ^ 1'h1;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T996;
  assign T996 = dmem_resp_valid & dmem_resp_fpu;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_ptw_status_ie = csr_io_status_ie;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_ie1 = csr_io_status_ie1;
  assign io_ptw_status_prv1 = csr_io_status_prv1;
  assign io_ptw_status_ie2 = csr_io_status_ie2;
  assign io_ptw_status_prv2 = csr_io_status_prv2;
  assign io_ptw_status_ie3 = csr_io_status_ie3;
  assign io_ptw_status_prv3 = csr_io_status_prv3;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_ptbr = csr_io_ptbr;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_dmem_req_bits_data = T997;
  assign T997 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_kill = T998;
  assign T998 = killm_common | mem_xcpt;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_tag = T1098;
  assign T1098 = {4'h0, T999};
  assign T999 = {ex_waddr, ex_ctrl_fp};
  assign io_dmem_req_bits_addr = T1000;
  assign T1000 = T1001;
  assign T1001 = {T1003, T1002};
  assign T1002 = alu_io_adder_out[6'h26:1'h0];
  assign T1003 = T1016 ? T1015 : T1004;
  assign T1004 = T1009 ? T1007 : T1005;
  assign T1005 = T1006[1'h0];
  assign T1006 = alu_io_adder_out[6'h27:6'h26];
  assign T1007 = T1008 == 2'h3;
  assign T1008 = T1006;
  assign T1009 = T1013 | T1010;
  assign T1010 = T1011 == 26'h3fffffe;
  assign T1011 = T1012;
  assign T1012 = ex_rs_0 >> 6'h26;
  assign T1013 = T1014 == 26'h3ffffff;
  assign T1014 = T1012;
  assign T1015 = T1006 != 2'h0;
  assign T1016 = T1018 | T1017;
  assign T1017 = T1012 == 26'h1;
  assign T1018 = T1012 == 26'h0;
  assign io_dmem_req_valid = T1019;
  assign T1019 = ex_reg_valid & ex_ctrl_mem;
  assign io_imem_invalidate = T1020;
  assign T1020 = wb_reg_valid & wb_ctrl_fence_i;
  assign T1021 = T650 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign T1022 = T649 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign T1023 = T65 ? id_ctrl_fence_i : ex_ctrl_fence_i;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_returnAddr = T1099;
  assign T1099 = mem_int_wdata[6'h26:1'h0];
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_isCall = T1024;
  assign T1024 = mem_ctrl_wxd & T1025;
  assign T1025 = mem_waddr[1'h0];
  assign io_imem_ras_update_valid = T1026;
  assign T1026 = T1028 & T1027;
  assign T1027 = take_pc_wb ^ 1'h1;
  assign T1028 = T1030 & T1029;
  assign T1029 = mem_npc_misaligned ^ 1'h1;
  assign T1030 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_pc = T1100;
  assign T1100 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_valid = T1031;
  assign T1031 = T1033 & T1032;
  assign T1032 = take_pc_wb ^ 1'h1;
  assign T1033 = mem_reg_valid & mem_ctrl_branch;
  assign io_imem_btb_update_bits_br_pc = T1101;
  assign T1101 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_isReturn = T1034;
  assign T1034 = mem_ctrl_jalr & T1035;
  assign T1035 = 5'h1 == T1036;
  assign T1036 = T1037 & 5'h19;
  assign T1037 = mem_reg_inst[5'h13:4'hf];
  assign io_imem_btb_update_bits_isJump = T1038;
  assign T1038 = mem_ctrl_jal | mem_ctrl_jalr;
  assign io_imem_btb_update_bits_target = T1102;
  assign T1102 = io_imem_req_bits_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_pc = T1103;
  assign T1103 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T1039 = T1042 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T1040 = T1041 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T1041 = T65 & io_imem_btb_resp_valid;
  assign T1042 = T649 & ex_reg_btb_hit;
  assign T1043 = T65 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T1044 = T1042 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T1045 = T1041 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T1046 = T1042 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T1047 = T1041 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T1048 = T1042 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T1049 = T1041 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign T1050 = T1042 ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign T1051 = T1041 ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign T1052 = T1042 ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign T1053 = T1041 ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T1054 = T1042 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T1055 = T1041 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T1056 = T649 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T1057;
  assign T1057 = T1059 & T1058;
  assign T1058 = take_pc_wb ^ 1'h1;
  assign T1059 = T1063 & T1060;
  assign T1060 = T1061 | mem_ctrl_jal;
  assign T1061 = T1062 | mem_ctrl_jalr;
  assign T1062 = mem_ctrl_branch & mem_br_taken;
  assign T1063 = T1064 & mem_wrong_npc;
  assign T1064 = mem_reg_valid & T1065;
  assign T1065 = mem_npc_misaligned ^ 1'h1;
  assign io_imem_resp_ready = T1066;
  assign T1066 = T1067 | csr_io_interrupt;
  assign T1067 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_bits_pc = T1068;
  assign T1068 = T1069;
  assign T1069 = T1071 ? csr_io_evec : T1070;
  assign T1070 = replay_wb ? wb_reg_pc : mem_npc;
  assign T1071 = wb_xcpt | csr_io_eret;
  assign io_imem_req_valid = take_pc;
  assign io_host_debug_stats_csr = csr_io_host_debug_stats_csr;
  assign io_host_csr_resp_bits = csr_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = csr_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = csr_io_host_csr_req_ready;
  CSRFile csr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( csr_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( csr_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( csr_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( csr_io_host_debug_stats_csr ),
       .io_rw_addr( T972 ),
       .io_rw_cmd( T971 ),
       .io_rw_rdata( csr_io_rw_rdata ),
       .io_rw_wdata( bypass_mux_2 ),
       .io_csr_stall( csr_io_csr_stall ),
       .io_csr_xcpt( csr_io_csr_xcpt ),
       .io_eret( csr_io_eret ),
       .io_status_sd( csr_io_status_sd ),
       .io_status_zero2( csr_io_status_zero2 ),
       .io_status_sd_rv32( csr_io_status_sd_rv32 ),
       .io_status_zero1( csr_io_status_zero1 ),
       .io_status_vm( csr_io_status_vm ),
       .io_status_mprv( csr_io_status_mprv ),
       .io_status_xs( csr_io_status_xs ),
       .io_status_fs( csr_io_status_fs ),
       .io_status_prv3( csr_io_status_prv3 ),
       .io_status_ie3( csr_io_status_ie3 ),
       .io_status_prv2( csr_io_status_prv2 ),
       .io_status_ie2( csr_io_status_ie2 ),
       .io_status_prv1( csr_io_status_prv1 ),
       .io_status_ie1( csr_io_status_ie1 ),
       .io_status_prv( csr_io_status_prv ),
       .io_status_ie( csr_io_status_ie ),
       .io_ptbr( csr_io_ptbr ),
       .io_evec( csr_io_evec ),
       .io_exception( wb_reg_xcpt ),
       .io_retire( wb_valid ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( wb_reg_cause ),
       .io_pc( wb_reg_pc ),
       .io_fatc( csr_io_fatc ),
       .io_time( csr_io_time ),
       .io_fcsr_rm( csr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_invalidate_lr( io_rocc_mem_invalidate_lr ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_autl_acquire_ready(  )
       .io_rocc_autl_acquire_valid( io_rocc_autl_acquire_valid ),
       .io_rocc_autl_acquire_bits_addr_block( io_rocc_autl_acquire_bits_addr_block ),
       .io_rocc_autl_acquire_bits_client_xact_id( io_rocc_autl_acquire_bits_client_xact_id ),
       .io_rocc_autl_acquire_bits_addr_beat( io_rocc_autl_acquire_bits_addr_beat ),
       .io_rocc_autl_acquire_bits_is_builtin_type( io_rocc_autl_acquire_bits_is_builtin_type ),
       .io_rocc_autl_acquire_bits_a_type( io_rocc_autl_acquire_bits_a_type ),
       .io_rocc_autl_acquire_bits_union( io_rocc_autl_acquire_bits_union ),
       .io_rocc_autl_acquire_bits_data( io_rocc_autl_acquire_bits_data ),
       .io_rocc_autl_grant_ready( io_rocc_autl_grant_ready ),
       //.io_rocc_autl_grant_valid(  )
       //.io_rocc_autl_grant_bits_addr_beat(  )
       //.io_rocc_autl_grant_bits_client_xact_id(  )
       //.io_rocc_autl_grant_bits_manager_xact_id(  )
       //.io_rocc_autl_grant_bits_is_builtin_type(  )
       //.io_rocc_autl_grant_bits_g_type(  )
       //.io_rocc_autl_grant_bits_data(  )
       //.io_rocc_fpu_req_ready(  )
       .io_rocc_fpu_req_valid( io_rocc_fpu_req_valid ),
       .io_rocc_fpu_req_bits_cmd( io_rocc_fpu_req_bits_cmd ),
       .io_rocc_fpu_req_bits_ldst( io_rocc_fpu_req_bits_ldst ),
       .io_rocc_fpu_req_bits_wen( io_rocc_fpu_req_bits_wen ),
       .io_rocc_fpu_req_bits_ren1( io_rocc_fpu_req_bits_ren1 ),
       .io_rocc_fpu_req_bits_ren2( io_rocc_fpu_req_bits_ren2 ),
       .io_rocc_fpu_req_bits_ren3( io_rocc_fpu_req_bits_ren3 ),
       .io_rocc_fpu_req_bits_swap12( io_rocc_fpu_req_bits_swap12 ),
       .io_rocc_fpu_req_bits_swap23( io_rocc_fpu_req_bits_swap23 ),
       .io_rocc_fpu_req_bits_single( io_rocc_fpu_req_bits_single ),
       .io_rocc_fpu_req_bits_fromint( io_rocc_fpu_req_bits_fromint ),
       .io_rocc_fpu_req_bits_toint( io_rocc_fpu_req_bits_toint ),
       .io_rocc_fpu_req_bits_fastpipe( io_rocc_fpu_req_bits_fastpipe ),
       .io_rocc_fpu_req_bits_fma( io_rocc_fpu_req_bits_fma ),
       .io_rocc_fpu_req_bits_div( io_rocc_fpu_req_bits_div ),
       .io_rocc_fpu_req_bits_sqrt( io_rocc_fpu_req_bits_sqrt ),
       .io_rocc_fpu_req_bits_round( io_rocc_fpu_req_bits_round ),
       .io_rocc_fpu_req_bits_wflags( io_rocc_fpu_req_bits_wflags ),
       .io_rocc_fpu_req_bits_rm( io_rocc_fpu_req_bits_rm ),
       .io_rocc_fpu_req_bits_typ( io_rocc_fpu_req_bits_typ ),
       .io_rocc_fpu_req_bits_in1( io_rocc_fpu_req_bits_in1 ),
       .io_rocc_fpu_req_bits_in2( io_rocc_fpu_req_bits_in2 ),
       .io_rocc_fpu_req_bits_in3( io_rocc_fpu_req_bits_in3 ),
       .io_rocc_fpu_resp_ready( io_rocc_fpu_resp_ready ),
       //.io_rocc_fpu_resp_valid(  )
       //.io_rocc_fpu_resp_bits_data(  )
       //.io_rocc_fpu_resp_bits_exc(  )
       //.io_rocc_exception(  )
       .io_rocc_csr_waddr( csr_io_rocc_csr_waddr ),
       .io_rocc_csr_wdata( csr_io_rocc_csr_wdata ),
       .io_rocc_csr_wen( csr_io_rocc_csr_wen ),
       //.io_rocc_host_id(  )
       .io_interrupt( csr_io_interrupt ),
       .io_interrupt_cause( csr_io_interrupt_cause )
  );
  ALU alu(
       .io_dw( ex_ctrl_alu_dw ),
       .io_fn( ex_ctrl_alu_fn ),
       .io_in2( T864 ),
       .io_in1( T834 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
       //.io_cmp_out(  )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( T833 ),
       .io_req_bits_fn( ex_ctrl_alu_fn ),
       .io_req_bits_dw( ex_ctrl_alu_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( ex_waddr ),
       .io_kill( T774 ),
       .io_resp_ready( T770 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );

  always @(posedge clk) begin
    if(T650) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T649) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data_0;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T48;
    end
    if(T650) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if(T649) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if(T65) begin
      ex_ctrl_rocc <= id_ctrl_rocc;
    end
    wb_reg_valid <= T66;
    if(T649) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    if(T65) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    mem_reg_valid <= T78;
    ex_reg_valid <= T80;
    if(T65) begin
      ex_reg_load_use <= id_load_use;
    end
    if(T649) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if(T65) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    if(T649) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if(T65) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if(T650) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if(T65) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if(T649) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if(T65) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if(T649) begin
      bypass_mux_1 <= alu_io_out;
    end
    if(T649) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if(T65) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if(T649) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T649) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if(T65) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if(T649) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if(T65) begin
      ex_reg_flush_pipe <= T243;
    end
    wb_reg_xcpt <= T262;
    mem_reg_xcpt <= T278;
    ex_reg_xcpt <= T281;
    ex_reg_xcpt_interrupt <= T412;
    mem_reg_xcpt_interrupt <= T416;
    wb_reg_replay <= T421;
    mem_reg_replay <= T424;
    if(reset) begin
      wb_reg_rocc_pending <= 1'h0;
    end else if(wb_reg_xcpt) begin
      wb_reg_rocc_pending <= 1'h0;
    end else if(wb_rocc_val) begin
      wb_reg_rocc_pending <= T441;
    end
    if(reset) begin
      R452 <= 32'h0;
    end else if(T489) begin
      R452 <= T485;
    end else if(T484) begin
      R452 <= T477;
    end else if(T459) begin
      R452 <= T456;
    end
    if(T650) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if(T649) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if(T65) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if(reset) begin
      R516 <= 32'h0;
    end else if(T527) begin
      R516 <= T519;
    end else if(ll_wen) begin
      R516 <= T503;
    end
    if(T650) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if(T650) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if(T649) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if(T649) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T65) begin
      ex_ctrl_mem_type <= id_ctrl_mem_type;
    end
    if(T65) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if(T649) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if(T65) begin
      ex_ctrl_csr <= id_csr;
    end else if(T65) begin
      ex_ctrl_csr <= id_ctrl_csr;
    end
    R654 <= R655;
    if(ex_reg_rs_bypass_1) begin
      R655 <= T708;
    end else begin
      R655 <= T656;
    end
    if(T697) begin
      ex_reg_rs_lsb_1 <= T671;
    end else if(T65) begin
      ex_reg_rs_lsb_1 <= T659;
    end
    if (T676)
      T674[T681] <= rf_wdata;
    if(T650) begin
      bypass_mux_2 <= T687;
    end
    if(T650) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if(T697) begin
      ex_reg_rs_msb_1 <= T707;
    end
    if(T65) begin
      ex_reg_rs_bypass_1 <= T700;
    end
    R719 <= R720;
    if(ex_reg_rs_bypass_0) begin
      R720 <= T749;
    end else begin
      R720 <= T721;
    end
    if(T739) begin
      ex_reg_rs_lsb_0 <= T732;
    end else if(T65) begin
      ex_reg_rs_lsb_0 <= T724;
    end
    if(T739) begin
      ex_reg_rs_msb_0 <= T748;
    end
    if(T65) begin
      ex_reg_rs_bypass_0 <= T742;
    end
    if(T650) begin
      wb_reg_pc <= mem_reg_pc;
    end
    R775 <= T776;
    if(T65) begin
      ex_ctrl_alu_dw <= id_ctrl_alu_dw;
    end
    if(T65) begin
      ex_ctrl_alu_fn <= id_ctrl_alu_fn;
    end
    if(T65) begin
      ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
    end
    if(T65) begin
      ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
    end
    if(T65) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(T985) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(T981) begin
      mem_reg_rs2 <= ex_rs_1;
    end
    if(T65) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if(T650) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if(T649) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if(T65) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if(T1042) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T1041) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(T65) begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T1042) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T1041) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T1042) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T1041) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T1042) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T1041) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T1042) begin
      mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
    end
    if(T1041) begin
      ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
    end
    if(T1042) begin
      mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
    end
    if(T1041) begin
      ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
    end
    if(T1042) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T1041) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T649) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T768, T766, T765, T763, T761, T760, T759, T757, T718, T716, T653, T652, T1);
// synthesis translate_on
`endif
  end
endmodule

module BTB(input clk, input reset,
    input  io_req_valid,
    input [38:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output io_resp_bits_mask,
    output io_resp_bits_bridx,
    output[38:0] io_resp_bits_target,
    output[5:0] io_resp_bits_entry,
    output[6:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_btb_update_valid,
    input  io_btb_update_bits_prediction_valid,
    input  io_btb_update_bits_prediction_bits_taken,
    input  io_btb_update_bits_prediction_bits_mask,
    input  io_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_btb_update_bits_prediction_bits_target,
    input [5:0] io_btb_update_bits_prediction_bits_entry,
    input [6:0] io_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_btb_update_bits_pc,
    input [38:0] io_btb_update_bits_target,
    input  io_btb_update_bits_taken,
    input  io_btb_update_bits_isJump,
    input  io_btb_update_bits_isReturn,
    input [38:0] io_btb_update_bits_br_pc,
    input  io_bht_update_valid,
    input  io_bht_update_bits_prediction_valid,
    input  io_bht_update_bits_prediction_bits_taken,
    input  io_bht_update_bits_prediction_bits_mask,
    input  io_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_bht_update_bits_prediction_bits_target,
    input [5:0] io_bht_update_bits_prediction_bits_entry,
    input [6:0] io_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_bht_update_bits_pc,
    input  io_bht_update_bits_taken,
    input  io_bht_update_bits_mispredict,
    input  io_ras_update_valid,
    input  io_ras_update_bits_isCall,
    input  io_ras_update_bits_isReturn,
    input [38:0] io_ras_update_bits_returnAddr,
    input  io_ras_update_bits_prediction_valid,
    input  io_ras_update_bits_prediction_bits_taken,
    input  io_ras_update_bits_prediction_bits_mask,
    input  io_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_ras_update_bits_prediction_bits_target,
    input [5:0] io_ras_update_bits_prediction_bits_entry,
    input [6:0] io_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_ras_update_bits_prediction_bits_bht_value,
    input  io_invalidate
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  reg [38:0] R4;
  wire[38:0] T5;
  wire T6;
  reg  R7;
  wire T2288;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10 [127:0];
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  reg [6:0] R25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[5:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg  isJump_61;
  wire T35;
  reg  R36;
  wire T37;
  wire T38;
  wire T39;
  wire[63:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  reg [5:0] nextRepl;
  wire[5:0] T2289;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire T46;
  wire T47;
  wire T48;
  reg [5:0] R49;
  wire[5:0] T50;
  reg  updateHit;
  wire T51;
  wire T52;
  wire[61:0] hits;
  wire[61:0] T53;
  wire[61:0] T54;
  wire[30:0] T55;
  wire[15:0] T56;
  wire[7:0] T57;
  wire[3:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[5:0] T61;
  wire[5:0] pageHit;
  reg [5:0] pageValid;
  wire[5:0] T2290;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] pageReplEn;
  wire[5:0] tgtPageReplEn;
  wire[5:0] tgtPageRepl;
  wire[5:0] T65;
  wire[5:0] T2291;
  wire T66;
  wire[5:0] T67;
  wire[4:0] T68;
  wire[5:0] idxPageUpdateOH;
  wire[5:0] idxPageRepl;
  wire[5:0] T2292;
  wire[7:0] T69;
  reg [2:0] R70;
  wire[2:0] T2293;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire[5:0] updatePageHit;
  wire[5:0] T76;
  wire[5:0] T77;
  wire[2:0] T78;
  wire[1:0] T79;
  wire T80;
  wire[26:0] T81;
  reg [38:0] R82;
  wire[38:0] T83;
  wire[26:0] T84;
  reg [26:0] pages [5:0];
  wire[26:0] T85;
  wire[26:0] T86;
  wire[26:0] T87;
  wire[26:0] T88;
  wire T89;
  wire[5:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire[26:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[26:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[26:0] T103;
  wire[26:0] T104;
  wire[26:0] T105;
  wire[26:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[26:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[26:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[26:0] T120;
  wire T121;
  wire[26:0] T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[26:0] T126;
  wire T127;
  wire[26:0] T128;
  wire T129;
  wire[26:0] T130;
  wire useUpdatePageHit;
  wire samePage;
  wire[26:0] T131;
  wire[26:0] T132;
  wire doTgtPageRepl;
  wire T133;
  wire usePageHit;
  wire[5:0] T134;
  wire[5:0] T135;
  wire T136;
  wire[5:0] idxPageReplEn;
  wire T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[2:0] T140;
  wire[1:0] T141;
  wire T142;
  wire[26:0] T143;
  wire[26:0] T144;
  wire T145;
  wire[26:0] T146;
  wire T147;
  wire[26:0] T148;
  wire[2:0] T149;
  wire[1:0] T150;
  wire T151;
  wire[26:0] T152;
  wire T153;
  wire[26:0] T154;
  wire T155;
  wire[26:0] T156;
  wire[5:0] idxPagesOH_0;
  wire[7:0] T157;
  wire[2:0] T158;
  reg [2:0] idxPages [61:0];
  wire[2:0] T159;
  wire[2:0] T2294;
  wire[1:0] T2295;
  wire T2296;
  wire[1:0] T2297;
  wire[1:0] T2298;
  wire[3:0] T2299;
  wire[3:0] T2300;
  wire[1:0] T2301;
  wire[1:0] T2302;
  wire T2303;
  wire T2304;
  wire T160;
  wire T161;
  wire T162;
  wire[5:0] T163;
  wire[5:0] idxPagesOH_1;
  wire[7:0] T164;
  wire[2:0] T165;
  wire[1:0] T166;
  wire T167;
  wire[5:0] T168;
  wire[5:0] idxPagesOH_2;
  wire[7:0] T169;
  wire[2:0] T170;
  wire T171;
  wire[5:0] T172;
  wire[5:0] idxPagesOH_3;
  wire[7:0] T173;
  wire[2:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire T177;
  wire[5:0] T178;
  wire[5:0] idxPagesOH_4;
  wire[7:0] T179;
  wire[2:0] T180;
  wire T181;
  wire[5:0] T182;
  wire[5:0] idxPagesOH_5;
  wire[7:0] T183;
  wire[2:0] T184;
  wire[1:0] T185;
  wire T186;
  wire[5:0] T187;
  wire[5:0] idxPagesOH_6;
  wire[7:0] T188;
  wire[2:0] T189;
  wire T190;
  wire[5:0] T191;
  wire[5:0] idxPagesOH_7;
  wire[7:0] T192;
  wire[2:0] T193;
  wire[7:0] T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire T197;
  wire[5:0] T198;
  wire[5:0] idxPagesOH_8;
  wire[7:0] T199;
  wire[2:0] T200;
  wire T201;
  wire[5:0] T202;
  wire[5:0] idxPagesOH_9;
  wire[7:0] T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[5:0] T207;
  wire[5:0] idxPagesOH_10;
  wire[7:0] T208;
  wire[2:0] T209;
  wire T210;
  wire[5:0] T211;
  wire[5:0] idxPagesOH_11;
  wire[7:0] T212;
  wire[2:0] T213;
  wire[3:0] T214;
  wire[1:0] T215;
  wire T216;
  wire[5:0] T217;
  wire[5:0] idxPagesOH_12;
  wire[7:0] T218;
  wire[2:0] T219;
  wire T220;
  wire[5:0] T221;
  wire[5:0] idxPagesOH_13;
  wire[7:0] T222;
  wire[2:0] T223;
  wire[1:0] T224;
  wire T225;
  wire[5:0] T226;
  wire[5:0] idxPagesOH_14;
  wire[7:0] T227;
  wire[2:0] T228;
  wire T229;
  wire[5:0] T230;
  wire[5:0] idxPagesOH_15;
  wire[7:0] T231;
  wire[2:0] T232;
  wire[14:0] T233;
  wire[7:0] T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire[5:0] T238;
  wire[5:0] idxPagesOH_16;
  wire[7:0] T239;
  wire[2:0] T240;
  wire T241;
  wire[5:0] T242;
  wire[5:0] idxPagesOH_17;
  wire[7:0] T243;
  wire[2:0] T244;
  wire[1:0] T245;
  wire T246;
  wire[5:0] T247;
  wire[5:0] idxPagesOH_18;
  wire[7:0] T248;
  wire[2:0] T249;
  wire T250;
  wire[5:0] T251;
  wire[5:0] idxPagesOH_19;
  wire[7:0] T252;
  wire[2:0] T253;
  wire[3:0] T254;
  wire[1:0] T255;
  wire T256;
  wire[5:0] T257;
  wire[5:0] idxPagesOH_20;
  wire[7:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[5:0] T261;
  wire[5:0] idxPagesOH_21;
  wire[7:0] T262;
  wire[2:0] T263;
  wire[1:0] T264;
  wire T265;
  wire[5:0] T266;
  wire[5:0] idxPagesOH_22;
  wire[7:0] T267;
  wire[2:0] T268;
  wire T269;
  wire[5:0] T270;
  wire[5:0] idxPagesOH_23;
  wire[7:0] T271;
  wire[2:0] T272;
  wire[6:0] T273;
  wire[3:0] T274;
  wire[1:0] T275;
  wire T276;
  wire[5:0] T277;
  wire[5:0] idxPagesOH_24;
  wire[7:0] T278;
  wire[2:0] T279;
  wire T280;
  wire[5:0] T281;
  wire[5:0] idxPagesOH_25;
  wire[7:0] T282;
  wire[2:0] T283;
  wire[1:0] T284;
  wire T285;
  wire[5:0] T286;
  wire[5:0] idxPagesOH_26;
  wire[7:0] T287;
  wire[2:0] T288;
  wire T289;
  wire[5:0] T290;
  wire[5:0] idxPagesOH_27;
  wire[7:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire[1:0] T294;
  wire T295;
  wire[5:0] T296;
  wire[5:0] idxPagesOH_28;
  wire[7:0] T297;
  wire[2:0] T298;
  wire T299;
  wire[5:0] T300;
  wire[5:0] idxPagesOH_29;
  wire[7:0] T301;
  wire[2:0] T302;
  wire T303;
  wire[5:0] T304;
  wire[5:0] idxPagesOH_30;
  wire[7:0] T305;
  wire[2:0] T306;
  wire[30:0] T307;
  wire[15:0] T308;
  wire[7:0] T309;
  wire[3:0] T310;
  wire[1:0] T311;
  wire T312;
  wire[5:0] T313;
  wire[5:0] idxPagesOH_31;
  wire[7:0] T314;
  wire[2:0] T315;
  wire T316;
  wire[5:0] T317;
  wire[5:0] idxPagesOH_32;
  wire[7:0] T318;
  wire[2:0] T319;
  wire[1:0] T320;
  wire T321;
  wire[5:0] T322;
  wire[5:0] idxPagesOH_33;
  wire[7:0] T323;
  wire[2:0] T324;
  wire T325;
  wire[5:0] T326;
  wire[5:0] idxPagesOH_34;
  wire[7:0] T327;
  wire[2:0] T328;
  wire[3:0] T329;
  wire[1:0] T330;
  wire T331;
  wire[5:0] T332;
  wire[5:0] idxPagesOH_35;
  wire[7:0] T333;
  wire[2:0] T334;
  wire T335;
  wire[5:0] T336;
  wire[5:0] idxPagesOH_36;
  wire[7:0] T337;
  wire[2:0] T338;
  wire[1:0] T339;
  wire T340;
  wire[5:0] T341;
  wire[5:0] idxPagesOH_37;
  wire[7:0] T342;
  wire[2:0] T343;
  wire T344;
  wire[5:0] T345;
  wire[5:0] idxPagesOH_38;
  wire[7:0] T346;
  wire[2:0] T347;
  wire[7:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire[5:0] T352;
  wire[5:0] idxPagesOH_39;
  wire[7:0] T353;
  wire[2:0] T354;
  wire T355;
  wire[5:0] T356;
  wire[5:0] idxPagesOH_40;
  wire[7:0] T357;
  wire[2:0] T358;
  wire[1:0] T359;
  wire T360;
  wire[5:0] T361;
  wire[5:0] idxPagesOH_41;
  wire[7:0] T362;
  wire[2:0] T363;
  wire T364;
  wire[5:0] T365;
  wire[5:0] idxPagesOH_42;
  wire[7:0] T366;
  wire[2:0] T367;
  wire[3:0] T368;
  wire[1:0] T369;
  wire T370;
  wire[5:0] T371;
  wire[5:0] idxPagesOH_43;
  wire[7:0] T372;
  wire[2:0] T373;
  wire T374;
  wire[5:0] T375;
  wire[5:0] idxPagesOH_44;
  wire[7:0] T376;
  wire[2:0] T377;
  wire[1:0] T378;
  wire T379;
  wire[5:0] T380;
  wire[5:0] idxPagesOH_45;
  wire[7:0] T381;
  wire[2:0] T382;
  wire T383;
  wire[5:0] T384;
  wire[5:0] idxPagesOH_46;
  wire[7:0] T385;
  wire[2:0] T386;
  wire[14:0] T387;
  wire[7:0] T388;
  wire[3:0] T389;
  wire[1:0] T390;
  wire T391;
  wire[5:0] T392;
  wire[5:0] idxPagesOH_47;
  wire[7:0] T393;
  wire[2:0] T394;
  wire T395;
  wire[5:0] T396;
  wire[5:0] idxPagesOH_48;
  wire[7:0] T397;
  wire[2:0] T398;
  wire[1:0] T399;
  wire T400;
  wire[5:0] T401;
  wire[5:0] idxPagesOH_49;
  wire[7:0] T402;
  wire[2:0] T403;
  wire T404;
  wire[5:0] T405;
  wire[5:0] idxPagesOH_50;
  wire[7:0] T406;
  wire[2:0] T407;
  wire[3:0] T408;
  wire[1:0] T409;
  wire T410;
  wire[5:0] T411;
  wire[5:0] idxPagesOH_51;
  wire[7:0] T412;
  wire[2:0] T413;
  wire T414;
  wire[5:0] T415;
  wire[5:0] idxPagesOH_52;
  wire[7:0] T416;
  wire[2:0] T417;
  wire[1:0] T418;
  wire T419;
  wire[5:0] T420;
  wire[5:0] idxPagesOH_53;
  wire[7:0] T421;
  wire[2:0] T422;
  wire T423;
  wire[5:0] T424;
  wire[5:0] idxPagesOH_54;
  wire[7:0] T425;
  wire[2:0] T426;
  wire[6:0] T427;
  wire[3:0] T428;
  wire[1:0] T429;
  wire T430;
  wire[5:0] T431;
  wire[5:0] idxPagesOH_55;
  wire[7:0] T432;
  wire[2:0] T433;
  wire T434;
  wire[5:0] T435;
  wire[5:0] idxPagesOH_56;
  wire[7:0] T436;
  wire[2:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[5:0] T440;
  wire[5:0] idxPagesOH_57;
  wire[7:0] T441;
  wire[2:0] T442;
  wire T443;
  wire[5:0] T444;
  wire[5:0] idxPagesOH_58;
  wire[7:0] T445;
  wire[2:0] T446;
  wire[2:0] T447;
  wire[1:0] T448;
  wire T449;
  wire[5:0] T450;
  wire[5:0] idxPagesOH_59;
  wire[7:0] T451;
  wire[2:0] T452;
  wire T453;
  wire[5:0] T454;
  wire[5:0] idxPagesOH_60;
  wire[7:0] T455;
  wire[2:0] T456;
  wire T457;
  wire[5:0] T458;
  wire[5:0] idxPagesOH_61;
  wire[7:0] T459;
  wire[2:0] T460;
  wire[61:0] T461;
  wire[61:0] T462;
  wire[61:0] T463;
  wire[30:0] T464;
  wire[15:0] T465;
  wire[7:0] T466;
  wire[3:0] T467;
  wire[1:0] T468;
  wire T469;
  wire[11:0] T470;
  wire[11:0] T471;
  reg [11:0] idxs [61:0];
  wire[11:0] T472;
  wire[11:0] T2305;
  wire T473;
  wire T474;
  wire T475;
  wire[11:0] T476;
  wire[1:0] T477;
  wire T478;
  wire[11:0] T479;
  wire T480;
  wire[11:0] T481;
  wire[3:0] T482;
  wire[1:0] T483;
  wire T484;
  wire[11:0] T485;
  wire T486;
  wire[11:0] T487;
  wire[1:0] T488;
  wire T489;
  wire[11:0] T490;
  wire T491;
  wire[11:0] T492;
  wire[7:0] T493;
  wire[3:0] T494;
  wire[1:0] T495;
  wire T496;
  wire[11:0] T497;
  wire T498;
  wire[11:0] T499;
  wire[1:0] T500;
  wire T501;
  wire[11:0] T502;
  wire T503;
  wire[11:0] T504;
  wire[3:0] T505;
  wire[1:0] T506;
  wire T507;
  wire[11:0] T508;
  wire T509;
  wire[11:0] T510;
  wire[1:0] T511;
  wire T512;
  wire[11:0] T513;
  wire T514;
  wire[11:0] T515;
  wire[14:0] T516;
  wire[7:0] T517;
  wire[3:0] T518;
  wire[1:0] T519;
  wire T520;
  wire[11:0] T521;
  wire T522;
  wire[11:0] T523;
  wire[1:0] T524;
  wire T525;
  wire[11:0] T526;
  wire T527;
  wire[11:0] T528;
  wire[3:0] T529;
  wire[1:0] T530;
  wire T531;
  wire[11:0] T532;
  wire T533;
  wire[11:0] T534;
  wire[1:0] T535;
  wire T536;
  wire[11:0] T537;
  wire T538;
  wire[11:0] T539;
  wire[6:0] T540;
  wire[3:0] T541;
  wire[1:0] T542;
  wire T543;
  wire[11:0] T544;
  wire T545;
  wire[11:0] T546;
  wire[1:0] T547;
  wire T548;
  wire[11:0] T549;
  wire T550;
  wire[11:0] T551;
  wire[2:0] T552;
  wire[1:0] T553;
  wire T554;
  wire[11:0] T555;
  wire T556;
  wire[11:0] T557;
  wire T558;
  wire[11:0] T559;
  wire[30:0] T560;
  wire[15:0] T561;
  wire[7:0] T562;
  wire[3:0] T563;
  wire[1:0] T564;
  wire T565;
  wire[11:0] T566;
  wire T567;
  wire[11:0] T568;
  wire[1:0] T569;
  wire T570;
  wire[11:0] T571;
  wire T572;
  wire[11:0] T573;
  wire[3:0] T574;
  wire[1:0] T575;
  wire T576;
  wire[11:0] T577;
  wire T578;
  wire[11:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[11:0] T582;
  wire T583;
  wire[11:0] T584;
  wire[7:0] T585;
  wire[3:0] T586;
  wire[1:0] T587;
  wire T588;
  wire[11:0] T589;
  wire T590;
  wire[11:0] T591;
  wire[1:0] T592;
  wire T593;
  wire[11:0] T594;
  wire T595;
  wire[11:0] T596;
  wire[3:0] T597;
  wire[1:0] T598;
  wire T599;
  wire[11:0] T600;
  wire T601;
  wire[11:0] T602;
  wire[1:0] T603;
  wire T604;
  wire[11:0] T605;
  wire T606;
  wire[11:0] T607;
  wire[14:0] T608;
  wire[7:0] T609;
  wire[3:0] T610;
  wire[1:0] T611;
  wire T612;
  wire[11:0] T613;
  wire T614;
  wire[11:0] T615;
  wire[1:0] T616;
  wire T617;
  wire[11:0] T618;
  wire T619;
  wire[11:0] T620;
  wire[3:0] T621;
  wire[1:0] T622;
  wire T623;
  wire[11:0] T624;
  wire T625;
  wire[11:0] T626;
  wire[1:0] T627;
  wire T628;
  wire[11:0] T629;
  wire T630;
  wire[11:0] T631;
  wire[6:0] T632;
  wire[3:0] T633;
  wire[1:0] T634;
  wire T635;
  wire[11:0] T636;
  wire T637;
  wire[11:0] T638;
  wire[1:0] T639;
  wire T640;
  wire[11:0] T641;
  wire T642;
  wire[11:0] T643;
  wire[2:0] T644;
  wire[1:0] T645;
  wire T646;
  wire[11:0] T647;
  wire T648;
  wire[11:0] T649;
  wire T650;
  wire[11:0] T651;
  reg [61:0] idxValid;
  wire[61:0] T2306;
  wire[63:0] T2307;
  wire[63:0] T652;
  wire[63:0] T653;
  wire[63:0] T2308;
  wire[63:0] T654;
  wire[63:0] T655;
  wire[63:0] T2309;
  wire[61:0] T656;
  wire[61:0] T657;
  wire[61:0] T658;
  wire[61:0] T659;
  wire[30:0] T660;
  wire[15:0] T661;
  wire[7:0] T662;
  wire[3:0] T663;
  wire[1:0] T664;
  wire T665;
  wire[5:0] T666;
  wire[5:0] T667;
  wire[5:0] tgtPagesOH_0;
  wire[7:0] T668;
  wire[2:0] T669;
  reg [2:0] tgtPages [61:0];
  wire[2:0] T670;
  wire[2:0] T2310;
  wire[1:0] T2311;
  wire T2312;
  wire[1:0] T2313;
  wire[1:0] T2314;
  wire[3:0] T2315;
  wire[3:0] T2316;
  wire[5:0] T671;
  wire[1:0] T2317;
  wire[1:0] T2318;
  wire T2319;
  wire T2320;
  wire T672;
  wire T673;
  wire T674;
  wire[5:0] T675;
  wire[5:0] T676;
  wire[5:0] tgtPagesOH_1;
  wire[7:0] T677;
  wire[2:0] T678;
  wire[1:0] T679;
  wire T680;
  wire[5:0] T681;
  wire[5:0] T682;
  wire[5:0] tgtPagesOH_2;
  wire[7:0] T683;
  wire[2:0] T684;
  wire T685;
  wire[5:0] T686;
  wire[5:0] T687;
  wire[5:0] tgtPagesOH_3;
  wire[7:0] T688;
  wire[2:0] T689;
  wire[3:0] T690;
  wire[1:0] T691;
  wire T692;
  wire[5:0] T693;
  wire[5:0] T694;
  wire[5:0] tgtPagesOH_4;
  wire[7:0] T695;
  wire[2:0] T696;
  wire T697;
  wire[5:0] T698;
  wire[5:0] T699;
  wire[5:0] tgtPagesOH_5;
  wire[7:0] T700;
  wire[2:0] T701;
  wire[1:0] T702;
  wire T703;
  wire[5:0] T704;
  wire[5:0] T705;
  wire[5:0] tgtPagesOH_6;
  wire[7:0] T706;
  wire[2:0] T707;
  wire T708;
  wire[5:0] T709;
  wire[5:0] T710;
  wire[5:0] tgtPagesOH_7;
  wire[7:0] T711;
  wire[2:0] T712;
  wire[7:0] T713;
  wire[3:0] T714;
  wire[1:0] T715;
  wire T716;
  wire[5:0] T717;
  wire[5:0] T718;
  wire[5:0] tgtPagesOH_8;
  wire[7:0] T719;
  wire[2:0] T720;
  wire T721;
  wire[5:0] T722;
  wire[5:0] T723;
  wire[5:0] tgtPagesOH_9;
  wire[7:0] T724;
  wire[2:0] T725;
  wire[1:0] T726;
  wire T727;
  wire[5:0] T728;
  wire[5:0] T729;
  wire[5:0] tgtPagesOH_10;
  wire[7:0] T730;
  wire[2:0] T731;
  wire T732;
  wire[5:0] T733;
  wire[5:0] T734;
  wire[5:0] tgtPagesOH_11;
  wire[7:0] T735;
  wire[2:0] T736;
  wire[3:0] T737;
  wire[1:0] T738;
  wire T739;
  wire[5:0] T740;
  wire[5:0] T741;
  wire[5:0] tgtPagesOH_12;
  wire[7:0] T742;
  wire[2:0] T743;
  wire T744;
  wire[5:0] T745;
  wire[5:0] T746;
  wire[5:0] tgtPagesOH_13;
  wire[7:0] T747;
  wire[2:0] T748;
  wire[1:0] T749;
  wire T750;
  wire[5:0] T751;
  wire[5:0] T752;
  wire[5:0] tgtPagesOH_14;
  wire[7:0] T753;
  wire[2:0] T754;
  wire T755;
  wire[5:0] T756;
  wire[5:0] T757;
  wire[5:0] tgtPagesOH_15;
  wire[7:0] T758;
  wire[2:0] T759;
  wire[14:0] T760;
  wire[7:0] T761;
  wire[3:0] T762;
  wire[1:0] T763;
  wire T764;
  wire[5:0] T765;
  wire[5:0] T766;
  wire[5:0] tgtPagesOH_16;
  wire[7:0] T767;
  wire[2:0] T768;
  wire T769;
  wire[5:0] T770;
  wire[5:0] T771;
  wire[5:0] tgtPagesOH_17;
  wire[7:0] T772;
  wire[2:0] T773;
  wire[1:0] T774;
  wire T775;
  wire[5:0] T776;
  wire[5:0] T777;
  wire[5:0] tgtPagesOH_18;
  wire[7:0] T778;
  wire[2:0] T779;
  wire T780;
  wire[5:0] T781;
  wire[5:0] T782;
  wire[5:0] tgtPagesOH_19;
  wire[7:0] T783;
  wire[2:0] T784;
  wire[3:0] T785;
  wire[1:0] T786;
  wire T787;
  wire[5:0] T788;
  wire[5:0] T789;
  wire[5:0] tgtPagesOH_20;
  wire[7:0] T790;
  wire[2:0] T791;
  wire T792;
  wire[5:0] T793;
  wire[5:0] T794;
  wire[5:0] tgtPagesOH_21;
  wire[7:0] T795;
  wire[2:0] T796;
  wire[1:0] T797;
  wire T798;
  wire[5:0] T799;
  wire[5:0] T800;
  wire[5:0] tgtPagesOH_22;
  wire[7:0] T801;
  wire[2:0] T802;
  wire T803;
  wire[5:0] T804;
  wire[5:0] T805;
  wire[5:0] tgtPagesOH_23;
  wire[7:0] T806;
  wire[2:0] T807;
  wire[6:0] T808;
  wire[3:0] T809;
  wire[1:0] T810;
  wire T811;
  wire[5:0] T812;
  wire[5:0] T813;
  wire[5:0] tgtPagesOH_24;
  wire[7:0] T814;
  wire[2:0] T815;
  wire T816;
  wire[5:0] T817;
  wire[5:0] T818;
  wire[5:0] tgtPagesOH_25;
  wire[7:0] T819;
  wire[2:0] T820;
  wire[1:0] T821;
  wire T822;
  wire[5:0] T823;
  wire[5:0] T824;
  wire[5:0] tgtPagesOH_26;
  wire[7:0] T825;
  wire[2:0] T826;
  wire T827;
  wire[5:0] T828;
  wire[5:0] T829;
  wire[5:0] tgtPagesOH_27;
  wire[7:0] T830;
  wire[2:0] T831;
  wire[2:0] T832;
  wire[1:0] T833;
  wire T834;
  wire[5:0] T835;
  wire[5:0] T836;
  wire[5:0] tgtPagesOH_28;
  wire[7:0] T837;
  wire[2:0] T838;
  wire T839;
  wire[5:0] T840;
  wire[5:0] T841;
  wire[5:0] tgtPagesOH_29;
  wire[7:0] T842;
  wire[2:0] T843;
  wire T844;
  wire[5:0] T845;
  wire[5:0] T846;
  wire[5:0] tgtPagesOH_30;
  wire[7:0] T847;
  wire[2:0] T848;
  wire[30:0] T849;
  wire[15:0] T850;
  wire[7:0] T851;
  wire[3:0] T852;
  wire[1:0] T853;
  wire T854;
  wire[5:0] T855;
  wire[5:0] T856;
  wire[5:0] tgtPagesOH_31;
  wire[7:0] T857;
  wire[2:0] T858;
  wire T859;
  wire[5:0] T860;
  wire[5:0] T861;
  wire[5:0] tgtPagesOH_32;
  wire[7:0] T862;
  wire[2:0] T863;
  wire[1:0] T864;
  wire T865;
  wire[5:0] T866;
  wire[5:0] T867;
  wire[5:0] tgtPagesOH_33;
  wire[7:0] T868;
  wire[2:0] T869;
  wire T870;
  wire[5:0] T871;
  wire[5:0] T872;
  wire[5:0] tgtPagesOH_34;
  wire[7:0] T873;
  wire[2:0] T874;
  wire[3:0] T875;
  wire[1:0] T876;
  wire T877;
  wire[5:0] T878;
  wire[5:0] T879;
  wire[5:0] tgtPagesOH_35;
  wire[7:0] T880;
  wire[2:0] T881;
  wire T882;
  wire[5:0] T883;
  wire[5:0] T884;
  wire[5:0] tgtPagesOH_36;
  wire[7:0] T885;
  wire[2:0] T886;
  wire[1:0] T887;
  wire T888;
  wire[5:0] T889;
  wire[5:0] T890;
  wire[5:0] tgtPagesOH_37;
  wire[7:0] T891;
  wire[2:0] T892;
  wire T893;
  wire[5:0] T894;
  wire[5:0] T895;
  wire[5:0] tgtPagesOH_38;
  wire[7:0] T896;
  wire[2:0] T897;
  wire[7:0] T898;
  wire[3:0] T899;
  wire[1:0] T900;
  wire T901;
  wire[5:0] T902;
  wire[5:0] T903;
  wire[5:0] tgtPagesOH_39;
  wire[7:0] T904;
  wire[2:0] T905;
  wire T906;
  wire[5:0] T907;
  wire[5:0] T908;
  wire[5:0] tgtPagesOH_40;
  wire[7:0] T909;
  wire[2:0] T910;
  wire[1:0] T911;
  wire T912;
  wire[5:0] T913;
  wire[5:0] T914;
  wire[5:0] tgtPagesOH_41;
  wire[7:0] T915;
  wire[2:0] T916;
  wire T917;
  wire[5:0] T918;
  wire[5:0] T919;
  wire[5:0] tgtPagesOH_42;
  wire[7:0] T920;
  wire[2:0] T921;
  wire[3:0] T922;
  wire[1:0] T923;
  wire T924;
  wire[5:0] T925;
  wire[5:0] T926;
  wire[5:0] tgtPagesOH_43;
  wire[7:0] T927;
  wire[2:0] T928;
  wire T929;
  wire[5:0] T930;
  wire[5:0] T931;
  wire[5:0] tgtPagesOH_44;
  wire[7:0] T932;
  wire[2:0] T933;
  wire[1:0] T934;
  wire T935;
  wire[5:0] T936;
  wire[5:0] T937;
  wire[5:0] tgtPagesOH_45;
  wire[7:0] T938;
  wire[2:0] T939;
  wire T940;
  wire[5:0] T941;
  wire[5:0] T942;
  wire[5:0] tgtPagesOH_46;
  wire[7:0] T943;
  wire[2:0] T944;
  wire[14:0] T945;
  wire[7:0] T946;
  wire[3:0] T947;
  wire[1:0] T948;
  wire T949;
  wire[5:0] T950;
  wire[5:0] T951;
  wire[5:0] tgtPagesOH_47;
  wire[7:0] T952;
  wire[2:0] T953;
  wire T954;
  wire[5:0] T955;
  wire[5:0] T956;
  wire[5:0] tgtPagesOH_48;
  wire[7:0] T957;
  wire[2:0] T958;
  wire[1:0] T959;
  wire T960;
  wire[5:0] T961;
  wire[5:0] T962;
  wire[5:0] tgtPagesOH_49;
  wire[7:0] T963;
  wire[2:0] T964;
  wire T965;
  wire[5:0] T966;
  wire[5:0] T967;
  wire[5:0] tgtPagesOH_50;
  wire[7:0] T968;
  wire[2:0] T969;
  wire[3:0] T970;
  wire[1:0] T971;
  wire T972;
  wire[5:0] T973;
  wire[5:0] T974;
  wire[5:0] tgtPagesOH_51;
  wire[7:0] T975;
  wire[2:0] T976;
  wire T977;
  wire[5:0] T978;
  wire[5:0] T979;
  wire[5:0] tgtPagesOH_52;
  wire[7:0] T980;
  wire[2:0] T981;
  wire[1:0] T982;
  wire T983;
  wire[5:0] T984;
  wire[5:0] T985;
  wire[5:0] tgtPagesOH_53;
  wire[7:0] T986;
  wire[2:0] T987;
  wire T988;
  wire[5:0] T989;
  wire[5:0] T990;
  wire[5:0] tgtPagesOH_54;
  wire[7:0] T991;
  wire[2:0] T992;
  wire[6:0] T993;
  wire[3:0] T994;
  wire[1:0] T995;
  wire T996;
  wire[5:0] T997;
  wire[5:0] T998;
  wire[5:0] tgtPagesOH_55;
  wire[7:0] T999;
  wire[2:0] T1000;
  wire T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[5:0] tgtPagesOH_56;
  wire[7:0] T1004;
  wire[2:0] T1005;
  wire[1:0] T1006;
  wire T1007;
  wire[5:0] T1008;
  wire[5:0] T1009;
  wire[5:0] tgtPagesOH_57;
  wire[7:0] T1010;
  wire[2:0] T1011;
  wire T1012;
  wire[5:0] T1013;
  wire[5:0] T1014;
  wire[5:0] tgtPagesOH_58;
  wire[7:0] T1015;
  wire[2:0] T1016;
  wire[2:0] T1017;
  wire[1:0] T1018;
  wire T1019;
  wire[5:0] T1020;
  wire[5:0] T1021;
  wire[5:0] tgtPagesOH_59;
  wire[7:0] T1022;
  wire[2:0] T1023;
  wire T1024;
  wire[5:0] T1025;
  wire[5:0] T1026;
  wire[5:0] tgtPagesOH_60;
  wire[7:0] T1027;
  wire[2:0] T1028;
  wire T1029;
  wire[5:0] T1030;
  wire[5:0] T1031;
  wire[5:0] tgtPagesOH_61;
  wire[7:0] T1032;
  wire[2:0] T1033;
  wire T1034;
  wire T1035;
  reg  isJump_60;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  reg  isJump_59;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  reg  isJump_58;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  reg  isJump_57;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  reg  isJump_56;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  reg  isJump_55;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  reg  isJump_54;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  reg  isJump_53;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  reg  isJump_52;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  reg  isJump_51;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  reg  isJump_50;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  reg  isJump_49;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  reg  isJump_48;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  reg  isJump_47;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  reg  isJump_46;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  reg  isJump_45;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  reg  isJump_44;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  reg  isJump_43;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  reg  isJump_42;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  reg  isJump_41;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  reg  isJump_40;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  reg  isJump_39;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  reg  isJump_38;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  reg  isJump_37;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  reg  isJump_36;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  reg  isJump_35;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  reg  isJump_34;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  reg  isJump_33;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  reg  isJump_32;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  reg  isJump_31;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  reg  isJump_30;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  reg  isJump_29;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  reg  isJump_28;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  reg  isJump_27;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  reg  isJump_26;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  reg  isJump_25;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  reg  isJump_24;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  reg  isJump_23;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  reg  isJump_22;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  reg  isJump_21;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  reg  isJump_20;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  reg  isJump_19;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  reg  isJump_18;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  reg  isJump_17;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  reg  isJump_16;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  reg  isJump_15;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  reg  isJump_14;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  reg  isJump_13;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  reg  isJump_12;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  reg  isJump_11;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  reg  isJump_10;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  reg  isJump_9;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  reg  isJump_8;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  reg  isJump_7;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  reg  isJump_6;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  reg  isJump_5;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  reg  isJump_4;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  reg  isJump_3;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  reg  isJump_2;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  reg  isJump_1;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  reg  isJump_0;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[6:0] T1400;
  wire[5:0] T1401;
  wire T1402;
  wire[6:0] T1403;
  wire[6:0] T1404;
  wire[5:0] T2321;
  wire[4:0] T2322;
  wire[3:0] T2323;
  wire[2:0] T2324;
  wire[1:0] T2325;
  wire T2326;
  wire[1:0] T2327;
  wire[1:0] T2328;
  wire[3:0] T2329;
  wire[3:0] T2330;
  wire[7:0] T2331;
  wire[7:0] T2332;
  wire[15:0] T2333;
  wire[15:0] T2334;
  wire[31:0] T2335;
  wire[31:0] T2336;
  wire[29:0] T2337;
  wire[15:0] T2338;
  wire[7:0] T2339;
  wire[3:0] T2340;
  wire[1:0] T2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  wire T2346;
  wire[38:0] T1406;
  wire[38:0] T1407;
  wire[38:0] T1408;
  wire[11:0] T1409;
  wire[11:0] T1410;
  wire[11:0] T1411;
  reg [11:0] tgts [61:0];
  wire[11:0] T1412;
  wire[11:0] T2347;
  wire T1413;
  wire T1414;
  wire T1415;
  wire[11:0] T1416;
  wire[11:0] T1417;
  wire[11:0] T1418;
  wire T1419;
  wire[11:0] T1420;
  wire[11:0] T1421;
  wire[11:0] T1422;
  wire T1423;
  wire[11:0] T1424;
  wire[11:0] T1425;
  wire[11:0] T1426;
  wire T1427;
  wire[11:0] T1428;
  wire[11:0] T1429;
  wire[11:0] T1430;
  wire T1431;
  wire[11:0] T1432;
  wire[11:0] T1433;
  wire[11:0] T1434;
  wire T1435;
  wire[11:0] T1436;
  wire[11:0] T1437;
  wire[11:0] T1438;
  wire T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[11:0] T1442;
  wire T1443;
  wire[11:0] T1444;
  wire[11:0] T1445;
  wire[11:0] T1446;
  wire T1447;
  wire[11:0] T1448;
  wire[11:0] T1449;
  wire[11:0] T1450;
  wire T1451;
  wire[11:0] T1452;
  wire[11:0] T1453;
  wire[11:0] T1454;
  wire T1455;
  wire[11:0] T1456;
  wire[11:0] T1457;
  wire[11:0] T1458;
  wire T1459;
  wire[11:0] T1460;
  wire[11:0] T1461;
  wire[11:0] T1462;
  wire T1463;
  wire[11:0] T1464;
  wire[11:0] T1465;
  wire[11:0] T1466;
  wire T1467;
  wire[11:0] T1468;
  wire[11:0] T1469;
  wire[11:0] T1470;
  wire T1471;
  wire[11:0] T1472;
  wire[11:0] T1473;
  wire[11:0] T1474;
  wire T1475;
  wire[11:0] T1476;
  wire[11:0] T1477;
  wire[11:0] T1478;
  wire T1479;
  wire[11:0] T1480;
  wire[11:0] T1481;
  wire[11:0] T1482;
  wire T1483;
  wire[11:0] T1484;
  wire[11:0] T1485;
  wire[11:0] T1486;
  wire T1487;
  wire[11:0] T1488;
  wire[11:0] T1489;
  wire[11:0] T1490;
  wire T1491;
  wire[11:0] T1492;
  wire[11:0] T1493;
  wire[11:0] T1494;
  wire T1495;
  wire[11:0] T1496;
  wire[11:0] T1497;
  wire[11:0] T1498;
  wire T1499;
  wire[11:0] T1500;
  wire[11:0] T1501;
  wire[11:0] T1502;
  wire T1503;
  wire[11:0] T1504;
  wire[11:0] T1505;
  wire[11:0] T1506;
  wire T1507;
  wire[11:0] T1508;
  wire[11:0] T1509;
  wire[11:0] T1510;
  wire T1511;
  wire[11:0] T1512;
  wire[11:0] T1513;
  wire[11:0] T1514;
  wire T1515;
  wire[11:0] T1516;
  wire[11:0] T1517;
  wire[11:0] T1518;
  wire T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[11:0] T1522;
  wire T1523;
  wire[11:0] T1524;
  wire[11:0] T1525;
  wire[11:0] T1526;
  wire T1527;
  wire[11:0] T1528;
  wire[11:0] T1529;
  wire[11:0] T1530;
  wire T1531;
  wire[11:0] T1532;
  wire[11:0] T1533;
  wire[11:0] T1534;
  wire T1535;
  wire[11:0] T1536;
  wire[11:0] T1537;
  wire[11:0] T1538;
  wire T1539;
  wire[11:0] T1540;
  wire[11:0] T1541;
  wire[11:0] T1542;
  wire T1543;
  wire[11:0] T1544;
  wire[11:0] T1545;
  wire[11:0] T1546;
  wire T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire[11:0] T1550;
  wire T1551;
  wire[11:0] T1552;
  wire[11:0] T1553;
  wire[11:0] T1554;
  wire T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire[11:0] T1558;
  wire T1559;
  wire[11:0] T1560;
  wire[11:0] T1561;
  wire[11:0] T1562;
  wire T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire[11:0] T1566;
  wire T1567;
  wire[11:0] T1568;
  wire[11:0] T1569;
  wire[11:0] T1570;
  wire T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire[11:0] T1574;
  wire T1575;
  wire[11:0] T1576;
  wire[11:0] T1577;
  wire[11:0] T1578;
  wire T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire[11:0] T1582;
  wire T1583;
  wire[11:0] T1584;
  wire[11:0] T1585;
  wire[11:0] T1586;
  wire T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire[11:0] T1590;
  wire T1591;
  wire[11:0] T1592;
  wire[11:0] T1593;
  wire[11:0] T1594;
  wire T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire[11:0] T1598;
  wire T1599;
  wire[11:0] T1600;
  wire[11:0] T1601;
  wire[11:0] T1602;
  wire T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire[11:0] T1606;
  wire T1607;
  wire[11:0] T1608;
  wire[11:0] T1609;
  wire[11:0] T1610;
  wire T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire[11:0] T1614;
  wire T1615;
  wire[11:0] T1616;
  wire[11:0] T1617;
  wire[11:0] T1618;
  wire T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire[11:0] T1622;
  wire T1623;
  wire[11:0] T1624;
  wire[11:0] T1625;
  wire[11:0] T1626;
  wire T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire[11:0] T1630;
  wire T1631;
  wire[11:0] T1632;
  wire[11:0] T1633;
  wire[11:0] T1634;
  wire T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire[11:0] T1638;
  wire T1639;
  wire[11:0] T1640;
  wire[11:0] T1641;
  wire[11:0] T1642;
  wire T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire[11:0] T1646;
  wire T1647;
  wire[11:0] T1648;
  wire[11:0] T1649;
  wire[11:0] T1650;
  wire T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire[11:0] T1654;
  wire T1655;
  wire[11:0] T1656;
  wire[11:0] T1657;
  wire T1658;
  wire[26:0] T1659;
  wire[26:0] T1660;
  wire[26:0] T1661;
  wire T1662;
  wire[5:0] T1663;
  wire[5:0] T1664;
  wire T1665;
  wire[5:0] T1666;
  wire[5:0] T1667;
  wire T1668;
  wire[5:0] T1669;
  wire[5:0] T1670;
  wire T1671;
  wire[5:0] T1672;
  wire[5:0] T1673;
  wire T1674;
  wire[5:0] T1675;
  wire[5:0] T1676;
  wire T1677;
  wire[5:0] T1678;
  wire[5:0] T1679;
  wire T1680;
  wire[5:0] T1681;
  wire[5:0] T1682;
  wire T1683;
  wire[5:0] T1684;
  wire[5:0] T1685;
  wire T1686;
  wire[5:0] T1687;
  wire[5:0] T1688;
  wire T1689;
  wire[5:0] T1690;
  wire[5:0] T1691;
  wire T1692;
  wire[5:0] T1693;
  wire[5:0] T1694;
  wire T1695;
  wire[5:0] T1696;
  wire[5:0] T1697;
  wire T1698;
  wire[5:0] T1699;
  wire[5:0] T1700;
  wire T1701;
  wire[5:0] T1702;
  wire[5:0] T1703;
  wire T1704;
  wire[5:0] T1705;
  wire[5:0] T1706;
  wire T1707;
  wire[5:0] T1708;
  wire[5:0] T1709;
  wire T1710;
  wire[5:0] T1711;
  wire[5:0] T1712;
  wire T1713;
  wire[5:0] T1714;
  wire[5:0] T1715;
  wire T1716;
  wire[5:0] T1717;
  wire[5:0] T1718;
  wire T1719;
  wire[5:0] T1720;
  wire[5:0] T1721;
  wire T1722;
  wire[5:0] T1723;
  wire[5:0] T1724;
  wire T1725;
  wire[5:0] T1726;
  wire[5:0] T1727;
  wire T1728;
  wire[5:0] T1729;
  wire[5:0] T1730;
  wire T1731;
  wire[5:0] T1732;
  wire[5:0] T1733;
  wire T1734;
  wire[5:0] T1735;
  wire[5:0] T1736;
  wire T1737;
  wire[5:0] T1738;
  wire[5:0] T1739;
  wire T1740;
  wire[5:0] T1741;
  wire[5:0] T1742;
  wire T1743;
  wire[5:0] T1744;
  wire[5:0] T1745;
  wire T1746;
  wire[5:0] T1747;
  wire[5:0] T1748;
  wire T1749;
  wire[5:0] T1750;
  wire[5:0] T1751;
  wire T1752;
  wire[5:0] T1753;
  wire[5:0] T1754;
  wire T1755;
  wire[5:0] T1756;
  wire[5:0] T1757;
  wire T1758;
  wire[5:0] T1759;
  wire[5:0] T1760;
  wire T1761;
  wire[5:0] T1762;
  wire[5:0] T1763;
  wire T1764;
  wire[5:0] T1765;
  wire[5:0] T1766;
  wire T1767;
  wire[5:0] T1768;
  wire[5:0] T1769;
  wire T1770;
  wire[5:0] T1771;
  wire[5:0] T1772;
  wire T1773;
  wire[5:0] T1774;
  wire[5:0] T1775;
  wire T1776;
  wire[5:0] T1777;
  wire[5:0] T1778;
  wire T1779;
  wire[5:0] T1780;
  wire[5:0] T1781;
  wire T1782;
  wire[5:0] T1783;
  wire[5:0] T1784;
  wire T1785;
  wire[5:0] T1786;
  wire[5:0] T1787;
  wire T1788;
  wire[5:0] T1789;
  wire[5:0] T1790;
  wire T1791;
  wire[5:0] T1792;
  wire[5:0] T1793;
  wire T1794;
  wire[5:0] T1795;
  wire[5:0] T1796;
  wire T1797;
  wire[5:0] T1798;
  wire[5:0] T1799;
  wire T1800;
  wire[5:0] T1801;
  wire[5:0] T1802;
  wire T1803;
  wire[5:0] T1804;
  wire[5:0] T1805;
  wire T1806;
  wire[5:0] T1807;
  wire[5:0] T1808;
  wire T1809;
  wire[5:0] T1810;
  wire[5:0] T1811;
  wire T1812;
  wire[5:0] T1813;
  wire[5:0] T1814;
  wire T1815;
  wire[5:0] T1816;
  wire[5:0] T1817;
  wire T1818;
  wire[5:0] T1819;
  wire[5:0] T1820;
  wire T1821;
  wire[5:0] T1822;
  wire[5:0] T1823;
  wire T1824;
  wire[5:0] T1825;
  wire[5:0] T1826;
  wire T1827;
  wire[5:0] T1828;
  wire[5:0] T1829;
  wire T1830;
  wire[5:0] T1831;
  wire[5:0] T1832;
  wire T1833;
  wire[5:0] T1834;
  wire[5:0] T1835;
  wire T1836;
  wire[5:0] T1837;
  wire[5:0] T1838;
  wire T1839;
  wire[5:0] T1840;
  wire[5:0] T1841;
  wire T1842;
  wire[5:0] T1843;
  wire[5:0] T1844;
  wire T1845;
  wire[5:0] T1846;
  wire T1847;
  wire[26:0] T1848;
  wire[26:0] T1849;
  wire[26:0] T1850;
  wire T1851;
  wire[26:0] T1852;
  wire[26:0] T1853;
  wire[26:0] T1854;
  wire T1855;
  wire[26:0] T1856;
  wire[26:0] T1857;
  wire[26:0] T1858;
  wire T1859;
  wire[26:0] T1860;
  wire[26:0] T1861;
  wire[26:0] T1862;
  wire T1863;
  wire[26:0] T1864;
  wire[26:0] T1865;
  wire T1866;
  wire[38:0] T1867;
  reg [38:0] R1868;
  wire[38:0] T1869;
  wire T1870;
  wire T1871;
  wire[1:0] T1872;
  wire T1873;
  wire T1874;
  reg  R1875;
  wire T2348;
  wire T1876;
  wire T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  reg [1:0] R1882;
  wire[1:0] T2349;
  wire[1:0] T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire[1:0] T1886;
  wire T1887;
  wire T1888;
  wire[1:0] T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire T1894;
  reg [38:0] R1895;
  wire[38:0] T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  reg  useRAS_61;
  wire T1903;
  reg  R1904;
  wire T1905;
  wire T1906;
  wire T1907;
  wire[63:0] T1908;
  wire[5:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  reg  useRAS_60;
  wire T1913;
  wire T1914;
  wire T1915;
  wire T1916;
  wire T1917;
  wire T1918;
  reg  useRAS_59;
  wire T1919;
  wire T1920;
  wire T1921;
  wire T1922;
  wire T1923;
  wire T1924;
  reg  useRAS_58;
  wire T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  reg  useRAS_57;
  wire T1931;
  wire T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  reg  useRAS_56;
  wire T1937;
  wire T1938;
  wire T1939;
  wire T1940;
  wire T1941;
  wire T1942;
  reg  useRAS_55;
  wire T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire T1947;
  wire T1948;
  reg  useRAS_54;
  wire T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  reg  useRAS_53;
  wire T1955;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  reg  useRAS_52;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  reg  useRAS_51;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  reg  useRAS_50;
  wire T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  reg  useRAS_49;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  reg  useRAS_48;
  wire T1985;
  wire T1986;
  wire T1987;
  wire T1988;
  wire T1989;
  wire T1990;
  reg  useRAS_47;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire T1996;
  reg  useRAS_46;
  wire T1997;
  wire T1998;
  wire T1999;
  wire T2000;
  wire T2001;
  wire T2002;
  reg  useRAS_45;
  wire T2003;
  wire T2004;
  wire T2005;
  wire T2006;
  wire T2007;
  wire T2008;
  reg  useRAS_44;
  wire T2009;
  wire T2010;
  wire T2011;
  wire T2012;
  wire T2013;
  wire T2014;
  reg  useRAS_43;
  wire T2015;
  wire T2016;
  wire T2017;
  wire T2018;
  wire T2019;
  wire T2020;
  reg  useRAS_42;
  wire T2021;
  wire T2022;
  wire T2023;
  wire T2024;
  wire T2025;
  wire T2026;
  reg  useRAS_41;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire T2032;
  reg  useRAS_40;
  wire T2033;
  wire T2034;
  wire T2035;
  wire T2036;
  wire T2037;
  wire T2038;
  reg  useRAS_39;
  wire T2039;
  wire T2040;
  wire T2041;
  wire T2042;
  wire T2043;
  wire T2044;
  reg  useRAS_38;
  wire T2045;
  wire T2046;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  reg  useRAS_37;
  wire T2051;
  wire T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  reg  useRAS_36;
  wire T2057;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  reg  useRAS_35;
  wire T2063;
  wire T2064;
  wire T2065;
  wire T2066;
  wire T2067;
  wire T2068;
  reg  useRAS_34;
  wire T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire T2073;
  wire T2074;
  reg  useRAS_33;
  wire T2075;
  wire T2076;
  wire T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  reg  useRAS_32;
  wire T2081;
  wire T2082;
  wire T2083;
  wire T2084;
  wire T2085;
  wire T2086;
  reg  useRAS_31;
  wire T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  reg  useRAS_30;
  wire T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire T2097;
  wire T2098;
  reg  useRAS_29;
  wire T2099;
  wire T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  reg  useRAS_28;
  wire T2105;
  wire T2106;
  wire T2107;
  wire T2108;
  wire T2109;
  wire T2110;
  reg  useRAS_27;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire T2116;
  reg  useRAS_26;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire T2121;
  wire T2122;
  reg  useRAS_25;
  wire T2123;
  wire T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  reg  useRAS_24;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire T2134;
  reg  useRAS_23;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire T2139;
  wire T2140;
  reg  useRAS_22;
  wire T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire T2145;
  wire T2146;
  reg  useRAS_21;
  wire T2147;
  wire T2148;
  wire T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  reg  useRAS_20;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  reg  useRAS_19;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  reg  useRAS_18;
  wire T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire T2169;
  wire T2170;
  reg  useRAS_17;
  wire T2171;
  wire T2172;
  wire T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  reg  useRAS_16;
  wire T2177;
  wire T2178;
  wire T2179;
  wire T2180;
  wire T2181;
  wire T2182;
  reg  useRAS_15;
  wire T2183;
  wire T2184;
  wire T2185;
  wire T2186;
  wire T2187;
  wire T2188;
  reg  useRAS_14;
  wire T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire T2193;
  wire T2194;
  reg  useRAS_13;
  wire T2195;
  wire T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  reg  useRAS_12;
  wire T2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  wire T2206;
  reg  useRAS_11;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  wire T2211;
  wire T2212;
  reg  useRAS_10;
  wire T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire T2217;
  wire T2218;
  reg  useRAS_9;
  wire T2219;
  wire T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  reg  useRAS_8;
  wire T2225;
  wire T2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  reg  useRAS_7;
  wire T2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  wire T2236;
  reg  useRAS_6;
  wire T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire T2241;
  wire T2242;
  reg  useRAS_5;
  wire T2243;
  wire T2244;
  wire T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  reg  useRAS_4;
  wire T2249;
  wire T2250;
  wire T2251;
  wire T2252;
  wire T2253;
  wire T2254;
  reg  useRAS_3;
  wire T2255;
  wire T2256;
  wire T2257;
  wire T2258;
  wire T2259;
  wire T2260;
  reg  useRAS_2;
  wire T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire T2265;
  wire T2266;
  reg  useRAS_1;
  wire T2267;
  wire T2268;
  wire T2269;
  wire T2270;
  wire T2271;
  reg  useRAS_0;
  wire T2272;
  wire T2273;
  wire T2274;
  wire T2275;
  wire T2276;
  wire T2277;
  wire T2278;
  wire T2279;
  reg  brIdx [61:0];
  wire T2280;
  wire T2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  wire T2286;
  wire T2287;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R7 = {1{$random}};
    for (initvar = 0; initvar < 128; initvar = initvar+1)
      T10[initvar] = {1{$random}};
    R25 = {1{$random}};
    isJump_61 = {1{$random}};
    R36 = {1{$random}};
    nextRepl = {1{$random}};
    R49 = {1{$random}};
    updateHit = {1{$random}};
    pageValid = {1{$random}};
    R70 = {1{$random}};
    R82 = {2{$random}};
    for (initvar = 0; initvar < 6; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {2{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    isJump_60 = {1{$random}};
    isJump_59 = {1{$random}};
    isJump_58 = {1{$random}};
    isJump_57 = {1{$random}};
    isJump_56 = {1{$random}};
    isJump_55 = {1{$random}};
    isJump_54 = {1{$random}};
    isJump_53 = {1{$random}};
    isJump_52 = {1{$random}};
    isJump_51 = {1{$random}};
    isJump_50 = {1{$random}};
    isJump_49 = {1{$random}};
    isJump_48 = {1{$random}};
    isJump_47 = {1{$random}};
    isJump_46 = {1{$random}};
    isJump_45 = {1{$random}};
    isJump_44 = {1{$random}};
    isJump_43 = {1{$random}};
    isJump_42 = {1{$random}};
    isJump_41 = {1{$random}};
    isJump_40 = {1{$random}};
    isJump_39 = {1{$random}};
    isJump_38 = {1{$random}};
    isJump_37 = {1{$random}};
    isJump_36 = {1{$random}};
    isJump_35 = {1{$random}};
    isJump_34 = {1{$random}};
    isJump_33 = {1{$random}};
    isJump_32 = {1{$random}};
    isJump_31 = {1{$random}};
    isJump_30 = {1{$random}};
    isJump_29 = {1{$random}};
    isJump_28 = {1{$random}};
    isJump_27 = {1{$random}};
    isJump_26 = {1{$random}};
    isJump_25 = {1{$random}};
    isJump_24 = {1{$random}};
    isJump_23 = {1{$random}};
    isJump_22 = {1{$random}};
    isJump_21 = {1{$random}};
    isJump_20 = {1{$random}};
    isJump_19 = {1{$random}};
    isJump_18 = {1{$random}};
    isJump_17 = {1{$random}};
    isJump_16 = {1{$random}};
    isJump_15 = {1{$random}};
    isJump_14 = {1{$random}};
    isJump_13 = {1{$random}};
    isJump_12 = {1{$random}};
    isJump_11 = {1{$random}};
    isJump_10 = {1{$random}};
    isJump_9 = {1{$random}};
    isJump_8 = {1{$random}};
    isJump_7 = {1{$random}};
    isJump_6 = {1{$random}};
    isJump_5 = {1{$random}};
    isJump_4 = {1{$random}};
    isJump_3 = {1{$random}};
    isJump_2 = {1{$random}};
    isJump_1 = {1{$random}};
    isJump_0 = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R1868 = {2{$random}};
    R1875 = {1{$random}};
    R1882 = {1{$random}};
    R1895 = {2{$random}};
    useRAS_61 = {1{$random}};
    R1904 = {1{$random}};
    useRAS_60 = {1{$random}};
    useRAS_59 = {1{$random}};
    useRAS_58 = {1{$random}};
    useRAS_57 = {1{$random}};
    useRAS_56 = {1{$random}};
    useRAS_55 = {1{$random}};
    useRAS_54 = {1{$random}};
    useRAS_53 = {1{$random}};
    useRAS_52 = {1{$random}};
    useRAS_51 = {1{$random}};
    useRAS_50 = {1{$random}};
    useRAS_49 = {1{$random}};
    useRAS_48 = {1{$random}};
    useRAS_47 = {1{$random}};
    useRAS_46 = {1{$random}};
    useRAS_45 = {1{$random}};
    useRAS_44 = {1{$random}};
    useRAS_43 = {1{$random}};
    useRAS_42 = {1{$random}};
    useRAS_41 = {1{$random}};
    useRAS_40 = {1{$random}};
    useRAS_39 = {1{$random}};
    useRAS_38 = {1{$random}};
    useRAS_37 = {1{$random}};
    useRAS_36 = {1{$random}};
    useRAS_35 = {1{$random}};
    useRAS_34 = {1{$random}};
    useRAS_33 = {1{$random}};
    useRAS_32 = {1{$random}};
    useRAS_31 = {1{$random}};
    useRAS_30 = {1{$random}};
    useRAS_29 = {1{$random}};
    useRAS_28 = {1{$random}};
    useRAS_27 = {1{$random}};
    useRAS_26 = {1{$random}};
    useRAS_25 = {1{$random}};
    useRAS_24 = {1{$random}};
    useRAS_23 = {1{$random}};
    useRAS_22 = {1{$random}};
    useRAS_21 = {1{$random}};
    useRAS_20 = {1{$random}};
    useRAS_19 = {1{$random}};
    useRAS_18 = {1{$random}};
    useRAS_17 = {1{$random}};
    useRAS_16 = {1{$random}};
    useRAS_15 = {1{$random}};
    useRAS_14 = {1{$random}};
    useRAS_13 = {1{$random}};
    useRAS_12 = {1{$random}};
    useRAS_11 = {1{$random}};
    useRAS_10 = {1{$random}};
    useRAS_9 = {1{$random}};
    useRAS_8 = {1{$random}};
    useRAS_7 = {1{$random}};
    useRAS_6 = {1{$random}};
    useRAS_5 = {1{$random}};
    useRAS_4 = {1{$random}};
    useRAS_3 = {1{$random}};
    useRAS_2 = {1{$random}};
    useRAS_1 = {1{$random}};
    useRAS_0 = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      brIdx[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_btb_update_valid ? io_btb_update_bits_target : R4;
  assign T6 = R7 ^ 1'h1;
  assign T2288 = reset ? 1'h0 : io_btb_update_valid;
  assign io_resp_bits_bht_value = T8;
  assign T8 = T9;
  assign T9 = T10[T24];
  assign T12 = {io_bht_update_bits_taken, T13};
  assign T13 = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = T17 | T16;
  assign T16 = io_bht_update_bits_prediction_bits_bht_value[1'h0];
  assign T17 = io_bht_update_bits_prediction_bits_bht_value[1'h1];
  assign T18 = T20 & T19;
  assign T19 = io_bht_update_bits_prediction_bits_bht_value[1'h0];
  assign T20 = io_bht_update_bits_prediction_bits_bht_value[1'h1];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22 = T23 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T23 = io_bht_update_bits_pc[4'h8:2'h2];
  assign T24 = T1403 ^ R25;
  assign T26 = T1402 ? T1400 : T27;
  assign T27 = T31 ? T28 : R25;
  assign T28 = {T30, T29};
  assign T29 = R25[3'h6:1'h1];
  assign T30 = T8[1'h0];
  assign T31 = T1399 & T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T1034 | T34;
  assign T34 = T52 ? isJump_61 : 1'h0;
  assign T35 = T38 ? R36 : isJump_61;
  assign T37 = io_btb_update_valid ? io_btb_update_bits_isJump : R36;
  assign T38 = R7 & T39;
  assign T39 = T40[6'h3d];
  assign T40 = 1'h1 << T41;
  assign T41 = T42;
  assign T42 = updateHit ? R49 : nextRepl;
  assign T2289 = reset ? 6'h0 : T43;
  assign T43 = T47 ? T44 : nextRepl;
  assign T44 = T46 ? 6'h0 : T45;
  assign T45 = nextRepl + 6'h1;
  assign T46 = nextRepl == 6'h3d;
  assign T47 = R7 & T48;
  assign T48 = updateHit ^ 1'h1;
  assign T50 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : R49;
  assign T51 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : updateHit;
  assign T52 = hits[6'h3d];
  assign hits = T461 & T53;
  assign T53 = T54;
  assign T54 = {T307, T55};
  assign T55 = {T233, T56};
  assign T56 = {T194, T57};
  assign T57 = {T175, T58};
  assign T58 = {T166, T59};
  assign T59 = {T162, T60};
  assign T60 = T61 != 6'h0;
  assign T61 = idxPagesOH_0 & pageHit;
  assign pageHit = T138 & pageValid;
  assign T2290 = reset ? 6'h0 : T62;
  assign T62 = io_invalidate ? 6'h0 : T63;
  assign T63 = T137 ? T64 : pageValid;
  assign T64 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 6'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T65;
  assign T65 = T67 | T2291;
  assign T2291 = {5'h0, T66};
  assign T66 = idxPageUpdateOH[3'h5];
  assign T67 = T68 << 1'h1;
  assign T68 = idxPageUpdateOH[3'h4:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T2292;
  assign T2292 = T69[3'h5:1'h0];
  assign T69 = 1'h1 << R70;
  assign T2293 = reset ? 3'h0 : T71;
  assign T71 = T75 ? T72 : R70;
  assign T72 = T74 ? 3'h0 : T73;
  assign T73 = R70 + 3'h1;
  assign T74 = R70 == 3'h5;
  assign T75 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = useUpdatePageHit ^ 1'h1;
  assign updatePageHit = T76 & pageValid;
  assign T76 = T77;
  assign T77 = {T123, T78};
  assign T78 = {T121, T79};
  assign T79 = {T119, T80};
  assign T80 = T84 == T81;
  assign T81 = R82 >> 4'hc;
  assign T83 = io_btb_update_valid ? io_btb_update_bits_pc : R82;
  assign T84 = pages[3'h0];
  assign T86 = T89 ? T88 : T87;
  assign T87 = R82 >> 4'hc;
  assign T88 = io_req_bits_addr >> 4'hc;
  assign T89 = T90 != 6'h0;
  assign T90 = idxPageUpdateOH & 6'h15;
  assign T91 = R7 & T92;
  assign T92 = T94 & T93;
  assign T93 = pageReplEn[3'h5];
  assign T94 = T89 ? doTgtPageRepl : doIdxPageRepl;
  assign T96 = R7 & T97;
  assign T97 = T94 & T98;
  assign T98 = pageReplEn[2'h3];
  assign T100 = R7 & T101;
  assign T101 = T94 & T102;
  assign T102 = pageReplEn[1'h1];
  assign T104 = T89 ? T106 : T105;
  assign T105 = io_req_bits_addr >> 4'hc;
  assign T106 = R82 >> 4'hc;
  assign T107 = R7 & T108;
  assign T108 = T110 & T109;
  assign T109 = pageReplEn[3'h4];
  assign T110 = T89 ? doIdxPageRepl : doTgtPageRepl;
  assign T112 = R7 & T113;
  assign T113 = T110 & T114;
  assign T114 = pageReplEn[2'h2];
  assign T116 = R7 & T117;
  assign T117 = T110 & T118;
  assign T118 = pageReplEn[1'h0];
  assign T119 = T120 == T81;
  assign T120 = pages[3'h1];
  assign T121 = T122 == T81;
  assign T122 = pages[3'h2];
  assign T123 = {T129, T124};
  assign T124 = {T127, T125};
  assign T125 = T126 == T81;
  assign T126 = pages[3'h3];
  assign T127 = T128 == T81;
  assign T128 = pages[3'h4];
  assign T129 = T130 == T81;
  assign T130 = pages[3'h5];
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign samePage = T132 == T131;
  assign T131 = io_req_bits_addr >> 4'hc;
  assign T132 = R82 >> 4'hc;
  assign doTgtPageRepl = T136 & T133;
  assign T133 = usePageHit ^ 1'h1;
  assign usePageHit = T134 != 6'h0;
  assign T134 = pageHit & T135;
  assign T135 = ~ idxPageReplEn;
  assign T136 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 6'h0;
  assign T137 = R7 & doPageRepl;
  assign T138 = T139;
  assign T139 = {T149, T140};
  assign T140 = {T147, T141};
  assign T141 = {T145, T142};
  assign T142 = T144 == T143;
  assign T143 = io_req_bits_addr >> 4'hc;
  assign T144 = pages[3'h0];
  assign T145 = T146 == T143;
  assign T146 = pages[3'h1];
  assign T147 = T148 == T143;
  assign T148 = pages[3'h2];
  assign T149 = {T155, T150};
  assign T150 = {T153, T151};
  assign T151 = T152 == T143;
  assign T152 = pages[3'h3];
  assign T153 = T154 == T143;
  assign T154 = pages[3'h4];
  assign T155 = T156 == T143;
  assign T156 = pages[3'h5];
  assign idxPagesOH_0 = T157[3'h5:1'h0];
  assign T157 = 1'h1 << T158;
  assign T158 = idxPages[6'h0];
  assign T2294 = {T2304, T2295};
  assign T2295 = {T2303, T2296};
  assign T2296 = T2297[1'h1];
  assign T2297 = T2302 | T2298;
  assign T2298 = T2299[1'h1:1'h0];
  assign T2299 = T2301 | T2300;
  assign T2300 = idxPageUpdateOH[2'h3:1'h0];
  assign T2301 = idxPageUpdateOH[3'h5:3'h4];
  assign T2302 = T2299[2'h3:2'h2];
  assign T2303 = T2302 != 2'h0;
  assign T2304 = T2301 != 2'h0;
  assign T160 = R7 & T161;
  assign T161 = T42 < 6'h3e;
  assign T162 = T163 != 6'h0;
  assign T163 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T164[3'h5:1'h0];
  assign T164 = 1'h1 << T165;
  assign T165 = idxPages[6'h1];
  assign T166 = {T171, T167};
  assign T167 = T168 != 6'h0;
  assign T168 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T169[3'h5:1'h0];
  assign T169 = 1'h1 << T170;
  assign T170 = idxPages[6'h2];
  assign T171 = T172 != 6'h0;
  assign T172 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T173[3'h5:1'h0];
  assign T173 = 1'h1 << T174;
  assign T174 = idxPages[6'h3];
  assign T175 = {T185, T176};
  assign T176 = {T181, T177};
  assign T177 = T178 != 6'h0;
  assign T178 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T179[3'h5:1'h0];
  assign T179 = 1'h1 << T180;
  assign T180 = idxPages[6'h4];
  assign T181 = T182 != 6'h0;
  assign T182 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T183[3'h5:1'h0];
  assign T183 = 1'h1 << T184;
  assign T184 = idxPages[6'h5];
  assign T185 = {T190, T186};
  assign T186 = T187 != 6'h0;
  assign T187 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T188[3'h5:1'h0];
  assign T188 = 1'h1 << T189;
  assign T189 = idxPages[6'h6];
  assign T190 = T191 != 6'h0;
  assign T191 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T192[3'h5:1'h0];
  assign T192 = 1'h1 << T193;
  assign T193 = idxPages[6'h7];
  assign T194 = {T214, T195};
  assign T195 = {T205, T196};
  assign T196 = {T201, T197};
  assign T197 = T198 != 6'h0;
  assign T198 = idxPagesOH_8 & pageHit;
  assign idxPagesOH_8 = T199[3'h5:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[6'h8];
  assign T201 = T202 != 6'h0;
  assign T202 = idxPagesOH_9 & pageHit;
  assign idxPagesOH_9 = T203[3'h5:1'h0];
  assign T203 = 1'h1 << T204;
  assign T204 = idxPages[6'h9];
  assign T205 = {T210, T206};
  assign T206 = T207 != 6'h0;
  assign T207 = idxPagesOH_10 & pageHit;
  assign idxPagesOH_10 = T208[3'h5:1'h0];
  assign T208 = 1'h1 << T209;
  assign T209 = idxPages[6'ha];
  assign T210 = T211 != 6'h0;
  assign T211 = idxPagesOH_11 & pageHit;
  assign idxPagesOH_11 = T212[3'h5:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = idxPages[6'hb];
  assign T214 = {T224, T215};
  assign T215 = {T220, T216};
  assign T216 = T217 != 6'h0;
  assign T217 = idxPagesOH_12 & pageHit;
  assign idxPagesOH_12 = T218[3'h5:1'h0];
  assign T218 = 1'h1 << T219;
  assign T219 = idxPages[6'hc];
  assign T220 = T221 != 6'h0;
  assign T221 = idxPagesOH_13 & pageHit;
  assign idxPagesOH_13 = T222[3'h5:1'h0];
  assign T222 = 1'h1 << T223;
  assign T223 = idxPages[6'hd];
  assign T224 = {T229, T225};
  assign T225 = T226 != 6'h0;
  assign T226 = idxPagesOH_14 & pageHit;
  assign idxPagesOH_14 = T227[3'h5:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = idxPages[6'he];
  assign T229 = T230 != 6'h0;
  assign T230 = idxPagesOH_15 & pageHit;
  assign idxPagesOH_15 = T231[3'h5:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = idxPages[6'hf];
  assign T233 = {T273, T234};
  assign T234 = {T254, T235};
  assign T235 = {T245, T236};
  assign T236 = {T241, T237};
  assign T237 = T238 != 6'h0;
  assign T238 = idxPagesOH_16 & pageHit;
  assign idxPagesOH_16 = T239[3'h5:1'h0];
  assign T239 = 1'h1 << T240;
  assign T240 = idxPages[6'h10];
  assign T241 = T242 != 6'h0;
  assign T242 = idxPagesOH_17 & pageHit;
  assign idxPagesOH_17 = T243[3'h5:1'h0];
  assign T243 = 1'h1 << T244;
  assign T244 = idxPages[6'h11];
  assign T245 = {T250, T246};
  assign T246 = T247 != 6'h0;
  assign T247 = idxPagesOH_18 & pageHit;
  assign idxPagesOH_18 = T248[3'h5:1'h0];
  assign T248 = 1'h1 << T249;
  assign T249 = idxPages[6'h12];
  assign T250 = T251 != 6'h0;
  assign T251 = idxPagesOH_19 & pageHit;
  assign idxPagesOH_19 = T252[3'h5:1'h0];
  assign T252 = 1'h1 << T253;
  assign T253 = idxPages[6'h13];
  assign T254 = {T264, T255};
  assign T255 = {T260, T256};
  assign T256 = T257 != 6'h0;
  assign T257 = idxPagesOH_20 & pageHit;
  assign idxPagesOH_20 = T258[3'h5:1'h0];
  assign T258 = 1'h1 << T259;
  assign T259 = idxPages[6'h14];
  assign T260 = T261 != 6'h0;
  assign T261 = idxPagesOH_21 & pageHit;
  assign idxPagesOH_21 = T262[3'h5:1'h0];
  assign T262 = 1'h1 << T263;
  assign T263 = idxPages[6'h15];
  assign T264 = {T269, T265};
  assign T265 = T266 != 6'h0;
  assign T266 = idxPagesOH_22 & pageHit;
  assign idxPagesOH_22 = T267[3'h5:1'h0];
  assign T267 = 1'h1 << T268;
  assign T268 = idxPages[6'h16];
  assign T269 = T270 != 6'h0;
  assign T270 = idxPagesOH_23 & pageHit;
  assign idxPagesOH_23 = T271[3'h5:1'h0];
  assign T271 = 1'h1 << T272;
  assign T272 = idxPages[6'h17];
  assign T273 = {T293, T274};
  assign T274 = {T284, T275};
  assign T275 = {T280, T276};
  assign T276 = T277 != 6'h0;
  assign T277 = idxPagesOH_24 & pageHit;
  assign idxPagesOH_24 = T278[3'h5:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = idxPages[6'h18];
  assign T280 = T281 != 6'h0;
  assign T281 = idxPagesOH_25 & pageHit;
  assign idxPagesOH_25 = T282[3'h5:1'h0];
  assign T282 = 1'h1 << T283;
  assign T283 = idxPages[6'h19];
  assign T284 = {T289, T285};
  assign T285 = T286 != 6'h0;
  assign T286 = idxPagesOH_26 & pageHit;
  assign idxPagesOH_26 = T287[3'h5:1'h0];
  assign T287 = 1'h1 << T288;
  assign T288 = idxPages[6'h1a];
  assign T289 = T290 != 6'h0;
  assign T290 = idxPagesOH_27 & pageHit;
  assign idxPagesOH_27 = T291[3'h5:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = idxPages[6'h1b];
  assign T293 = {T303, T294};
  assign T294 = {T299, T295};
  assign T295 = T296 != 6'h0;
  assign T296 = idxPagesOH_28 & pageHit;
  assign idxPagesOH_28 = T297[3'h5:1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = idxPages[6'h1c];
  assign T299 = T300 != 6'h0;
  assign T300 = idxPagesOH_29 & pageHit;
  assign idxPagesOH_29 = T301[3'h5:1'h0];
  assign T301 = 1'h1 << T302;
  assign T302 = idxPages[6'h1d];
  assign T303 = T304 != 6'h0;
  assign T304 = idxPagesOH_30 & pageHit;
  assign idxPagesOH_30 = T305[3'h5:1'h0];
  assign T305 = 1'h1 << T306;
  assign T306 = idxPages[6'h1e];
  assign T307 = {T387, T308};
  assign T308 = {T348, T309};
  assign T309 = {T329, T310};
  assign T310 = {T320, T311};
  assign T311 = {T316, T312};
  assign T312 = T313 != 6'h0;
  assign T313 = idxPagesOH_31 & pageHit;
  assign idxPagesOH_31 = T314[3'h5:1'h0];
  assign T314 = 1'h1 << T315;
  assign T315 = idxPages[6'h1f];
  assign T316 = T317 != 6'h0;
  assign T317 = idxPagesOH_32 & pageHit;
  assign idxPagesOH_32 = T318[3'h5:1'h0];
  assign T318 = 1'h1 << T319;
  assign T319 = idxPages[6'h20];
  assign T320 = {T325, T321};
  assign T321 = T322 != 6'h0;
  assign T322 = idxPagesOH_33 & pageHit;
  assign idxPagesOH_33 = T323[3'h5:1'h0];
  assign T323 = 1'h1 << T324;
  assign T324 = idxPages[6'h21];
  assign T325 = T326 != 6'h0;
  assign T326 = idxPagesOH_34 & pageHit;
  assign idxPagesOH_34 = T327[3'h5:1'h0];
  assign T327 = 1'h1 << T328;
  assign T328 = idxPages[6'h22];
  assign T329 = {T339, T330};
  assign T330 = {T335, T331};
  assign T331 = T332 != 6'h0;
  assign T332 = idxPagesOH_35 & pageHit;
  assign idxPagesOH_35 = T333[3'h5:1'h0];
  assign T333 = 1'h1 << T334;
  assign T334 = idxPages[6'h23];
  assign T335 = T336 != 6'h0;
  assign T336 = idxPagesOH_36 & pageHit;
  assign idxPagesOH_36 = T337[3'h5:1'h0];
  assign T337 = 1'h1 << T338;
  assign T338 = idxPages[6'h24];
  assign T339 = {T344, T340};
  assign T340 = T341 != 6'h0;
  assign T341 = idxPagesOH_37 & pageHit;
  assign idxPagesOH_37 = T342[3'h5:1'h0];
  assign T342 = 1'h1 << T343;
  assign T343 = idxPages[6'h25];
  assign T344 = T345 != 6'h0;
  assign T345 = idxPagesOH_38 & pageHit;
  assign idxPagesOH_38 = T346[3'h5:1'h0];
  assign T346 = 1'h1 << T347;
  assign T347 = idxPages[6'h26];
  assign T348 = {T368, T349};
  assign T349 = {T359, T350};
  assign T350 = {T355, T351};
  assign T351 = T352 != 6'h0;
  assign T352 = idxPagesOH_39 & pageHit;
  assign idxPagesOH_39 = T353[3'h5:1'h0];
  assign T353 = 1'h1 << T354;
  assign T354 = idxPages[6'h27];
  assign T355 = T356 != 6'h0;
  assign T356 = idxPagesOH_40 & pageHit;
  assign idxPagesOH_40 = T357[3'h5:1'h0];
  assign T357 = 1'h1 << T358;
  assign T358 = idxPages[6'h28];
  assign T359 = {T364, T360};
  assign T360 = T361 != 6'h0;
  assign T361 = idxPagesOH_41 & pageHit;
  assign idxPagesOH_41 = T362[3'h5:1'h0];
  assign T362 = 1'h1 << T363;
  assign T363 = idxPages[6'h29];
  assign T364 = T365 != 6'h0;
  assign T365 = idxPagesOH_42 & pageHit;
  assign idxPagesOH_42 = T366[3'h5:1'h0];
  assign T366 = 1'h1 << T367;
  assign T367 = idxPages[6'h2a];
  assign T368 = {T378, T369};
  assign T369 = {T374, T370};
  assign T370 = T371 != 6'h0;
  assign T371 = idxPagesOH_43 & pageHit;
  assign idxPagesOH_43 = T372[3'h5:1'h0];
  assign T372 = 1'h1 << T373;
  assign T373 = idxPages[6'h2b];
  assign T374 = T375 != 6'h0;
  assign T375 = idxPagesOH_44 & pageHit;
  assign idxPagesOH_44 = T376[3'h5:1'h0];
  assign T376 = 1'h1 << T377;
  assign T377 = idxPages[6'h2c];
  assign T378 = {T383, T379};
  assign T379 = T380 != 6'h0;
  assign T380 = idxPagesOH_45 & pageHit;
  assign idxPagesOH_45 = T381[3'h5:1'h0];
  assign T381 = 1'h1 << T382;
  assign T382 = idxPages[6'h2d];
  assign T383 = T384 != 6'h0;
  assign T384 = idxPagesOH_46 & pageHit;
  assign idxPagesOH_46 = T385[3'h5:1'h0];
  assign T385 = 1'h1 << T386;
  assign T386 = idxPages[6'h2e];
  assign T387 = {T427, T388};
  assign T388 = {T408, T389};
  assign T389 = {T399, T390};
  assign T390 = {T395, T391};
  assign T391 = T392 != 6'h0;
  assign T392 = idxPagesOH_47 & pageHit;
  assign idxPagesOH_47 = T393[3'h5:1'h0];
  assign T393 = 1'h1 << T394;
  assign T394 = idxPages[6'h2f];
  assign T395 = T396 != 6'h0;
  assign T396 = idxPagesOH_48 & pageHit;
  assign idxPagesOH_48 = T397[3'h5:1'h0];
  assign T397 = 1'h1 << T398;
  assign T398 = idxPages[6'h30];
  assign T399 = {T404, T400};
  assign T400 = T401 != 6'h0;
  assign T401 = idxPagesOH_49 & pageHit;
  assign idxPagesOH_49 = T402[3'h5:1'h0];
  assign T402 = 1'h1 << T403;
  assign T403 = idxPages[6'h31];
  assign T404 = T405 != 6'h0;
  assign T405 = idxPagesOH_50 & pageHit;
  assign idxPagesOH_50 = T406[3'h5:1'h0];
  assign T406 = 1'h1 << T407;
  assign T407 = idxPages[6'h32];
  assign T408 = {T418, T409};
  assign T409 = {T414, T410};
  assign T410 = T411 != 6'h0;
  assign T411 = idxPagesOH_51 & pageHit;
  assign idxPagesOH_51 = T412[3'h5:1'h0];
  assign T412 = 1'h1 << T413;
  assign T413 = idxPages[6'h33];
  assign T414 = T415 != 6'h0;
  assign T415 = idxPagesOH_52 & pageHit;
  assign idxPagesOH_52 = T416[3'h5:1'h0];
  assign T416 = 1'h1 << T417;
  assign T417 = idxPages[6'h34];
  assign T418 = {T423, T419};
  assign T419 = T420 != 6'h0;
  assign T420 = idxPagesOH_53 & pageHit;
  assign idxPagesOH_53 = T421[3'h5:1'h0];
  assign T421 = 1'h1 << T422;
  assign T422 = idxPages[6'h35];
  assign T423 = T424 != 6'h0;
  assign T424 = idxPagesOH_54 & pageHit;
  assign idxPagesOH_54 = T425[3'h5:1'h0];
  assign T425 = 1'h1 << T426;
  assign T426 = idxPages[6'h36];
  assign T427 = {T447, T428};
  assign T428 = {T438, T429};
  assign T429 = {T434, T430};
  assign T430 = T431 != 6'h0;
  assign T431 = idxPagesOH_55 & pageHit;
  assign idxPagesOH_55 = T432[3'h5:1'h0];
  assign T432 = 1'h1 << T433;
  assign T433 = idxPages[6'h37];
  assign T434 = T435 != 6'h0;
  assign T435 = idxPagesOH_56 & pageHit;
  assign idxPagesOH_56 = T436[3'h5:1'h0];
  assign T436 = 1'h1 << T437;
  assign T437 = idxPages[6'h38];
  assign T438 = {T443, T439};
  assign T439 = T440 != 6'h0;
  assign T440 = idxPagesOH_57 & pageHit;
  assign idxPagesOH_57 = T441[3'h5:1'h0];
  assign T441 = 1'h1 << T442;
  assign T442 = idxPages[6'h39];
  assign T443 = T444 != 6'h0;
  assign T444 = idxPagesOH_58 & pageHit;
  assign idxPagesOH_58 = T445[3'h5:1'h0];
  assign T445 = 1'h1 << T446;
  assign T446 = idxPages[6'h3a];
  assign T447 = {T457, T448};
  assign T448 = {T453, T449};
  assign T449 = T450 != 6'h0;
  assign T450 = idxPagesOH_59 & pageHit;
  assign idxPagesOH_59 = T451[3'h5:1'h0];
  assign T451 = 1'h1 << T452;
  assign T452 = idxPages[6'h3b];
  assign T453 = T454 != 6'h0;
  assign T454 = idxPagesOH_60 & pageHit;
  assign idxPagesOH_60 = T455[3'h5:1'h0];
  assign T455 = 1'h1 << T456;
  assign T456 = idxPages[6'h3c];
  assign T457 = T458 != 6'h0;
  assign T458 = idxPagesOH_61 & pageHit;
  assign idxPagesOH_61 = T459[3'h5:1'h0];
  assign T459 = 1'h1 << T460;
  assign T460 = idxPages[6'h3d];
  assign T461 = idxValid & T462;
  assign T462 = T463;
  assign T463 = {T560, T464};
  assign T464 = {T516, T465};
  assign T465 = {T493, T466};
  assign T466 = {T482, T467};
  assign T467 = {T477, T468};
  assign T468 = {T475, T469};
  assign T469 = T471 == T470;
  assign T470 = io_req_bits_addr[4'hb:1'h0];
  assign T471 = idxs[6'h0];
  assign T2305 = R82[4'hb:1'h0];
  assign T473 = R7 & T474;
  assign T474 = T42 < 6'h3e;
  assign T475 = T476 == T470;
  assign T476 = idxs[6'h1];
  assign T477 = {T480, T478};
  assign T478 = T479 == T470;
  assign T479 = idxs[6'h2];
  assign T480 = T481 == T470;
  assign T481 = idxs[6'h3];
  assign T482 = {T488, T483};
  assign T483 = {T486, T484};
  assign T484 = T485 == T470;
  assign T485 = idxs[6'h4];
  assign T486 = T487 == T470;
  assign T487 = idxs[6'h5];
  assign T488 = {T491, T489};
  assign T489 = T490 == T470;
  assign T490 = idxs[6'h6];
  assign T491 = T492 == T470;
  assign T492 = idxs[6'h7];
  assign T493 = {T505, T494};
  assign T494 = {T500, T495};
  assign T495 = {T498, T496};
  assign T496 = T497 == T470;
  assign T497 = idxs[6'h8];
  assign T498 = T499 == T470;
  assign T499 = idxs[6'h9];
  assign T500 = {T503, T501};
  assign T501 = T502 == T470;
  assign T502 = idxs[6'ha];
  assign T503 = T504 == T470;
  assign T504 = idxs[6'hb];
  assign T505 = {T511, T506};
  assign T506 = {T509, T507};
  assign T507 = T508 == T470;
  assign T508 = idxs[6'hc];
  assign T509 = T510 == T470;
  assign T510 = idxs[6'hd];
  assign T511 = {T514, T512};
  assign T512 = T513 == T470;
  assign T513 = idxs[6'he];
  assign T514 = T515 == T470;
  assign T515 = idxs[6'hf];
  assign T516 = {T540, T517};
  assign T517 = {T529, T518};
  assign T518 = {T524, T519};
  assign T519 = {T522, T520};
  assign T520 = T521 == T470;
  assign T521 = idxs[6'h10];
  assign T522 = T523 == T470;
  assign T523 = idxs[6'h11];
  assign T524 = {T527, T525};
  assign T525 = T526 == T470;
  assign T526 = idxs[6'h12];
  assign T527 = T528 == T470;
  assign T528 = idxs[6'h13];
  assign T529 = {T535, T530};
  assign T530 = {T533, T531};
  assign T531 = T532 == T470;
  assign T532 = idxs[6'h14];
  assign T533 = T534 == T470;
  assign T534 = idxs[6'h15];
  assign T535 = {T538, T536};
  assign T536 = T537 == T470;
  assign T537 = idxs[6'h16];
  assign T538 = T539 == T470;
  assign T539 = idxs[6'h17];
  assign T540 = {T552, T541};
  assign T541 = {T547, T542};
  assign T542 = {T545, T543};
  assign T543 = T544 == T470;
  assign T544 = idxs[6'h18];
  assign T545 = T546 == T470;
  assign T546 = idxs[6'h19];
  assign T547 = {T550, T548};
  assign T548 = T549 == T470;
  assign T549 = idxs[6'h1a];
  assign T550 = T551 == T470;
  assign T551 = idxs[6'h1b];
  assign T552 = {T558, T553};
  assign T553 = {T556, T554};
  assign T554 = T555 == T470;
  assign T555 = idxs[6'h1c];
  assign T556 = T557 == T470;
  assign T557 = idxs[6'h1d];
  assign T558 = T559 == T470;
  assign T559 = idxs[6'h1e];
  assign T560 = {T608, T561};
  assign T561 = {T585, T562};
  assign T562 = {T574, T563};
  assign T563 = {T569, T564};
  assign T564 = {T567, T565};
  assign T565 = T566 == T470;
  assign T566 = idxs[6'h1f];
  assign T567 = T568 == T470;
  assign T568 = idxs[6'h20];
  assign T569 = {T572, T570};
  assign T570 = T571 == T470;
  assign T571 = idxs[6'h21];
  assign T572 = T573 == T470;
  assign T573 = idxs[6'h22];
  assign T574 = {T580, T575};
  assign T575 = {T578, T576};
  assign T576 = T577 == T470;
  assign T577 = idxs[6'h23];
  assign T578 = T579 == T470;
  assign T579 = idxs[6'h24];
  assign T580 = {T583, T581};
  assign T581 = T582 == T470;
  assign T582 = idxs[6'h25];
  assign T583 = T584 == T470;
  assign T584 = idxs[6'h26];
  assign T585 = {T597, T586};
  assign T586 = {T592, T587};
  assign T587 = {T590, T588};
  assign T588 = T589 == T470;
  assign T589 = idxs[6'h27];
  assign T590 = T591 == T470;
  assign T591 = idxs[6'h28];
  assign T592 = {T595, T593};
  assign T593 = T594 == T470;
  assign T594 = idxs[6'h29];
  assign T595 = T596 == T470;
  assign T596 = idxs[6'h2a];
  assign T597 = {T603, T598};
  assign T598 = {T601, T599};
  assign T599 = T600 == T470;
  assign T600 = idxs[6'h2b];
  assign T601 = T602 == T470;
  assign T602 = idxs[6'h2c];
  assign T603 = {T606, T604};
  assign T604 = T605 == T470;
  assign T605 = idxs[6'h2d];
  assign T606 = T607 == T470;
  assign T607 = idxs[6'h2e];
  assign T608 = {T632, T609};
  assign T609 = {T621, T610};
  assign T610 = {T616, T611};
  assign T611 = {T614, T612};
  assign T612 = T613 == T470;
  assign T613 = idxs[6'h2f];
  assign T614 = T615 == T470;
  assign T615 = idxs[6'h30];
  assign T616 = {T619, T617};
  assign T617 = T618 == T470;
  assign T618 = idxs[6'h31];
  assign T619 = T620 == T470;
  assign T620 = idxs[6'h32];
  assign T621 = {T627, T622};
  assign T622 = {T625, T623};
  assign T623 = T624 == T470;
  assign T624 = idxs[6'h33];
  assign T625 = T626 == T470;
  assign T626 = idxs[6'h34];
  assign T627 = {T630, T628};
  assign T628 = T629 == T470;
  assign T629 = idxs[6'h35];
  assign T630 = T631 == T470;
  assign T631 = idxs[6'h36];
  assign T632 = {T644, T633};
  assign T633 = {T639, T634};
  assign T634 = {T637, T635};
  assign T635 = T636 == T470;
  assign T636 = idxs[6'h37];
  assign T637 = T638 == T470;
  assign T638 = idxs[6'h38];
  assign T639 = {T642, T640};
  assign T640 = T641 == T470;
  assign T641 = idxs[6'h39];
  assign T642 = T643 == T470;
  assign T643 = idxs[6'h3a];
  assign T644 = {T650, T645};
  assign T645 = {T648, T646};
  assign T646 = T647 == T470;
  assign T647 = idxs[6'h3b];
  assign T648 = T649 == T470;
  assign T649 = idxs[6'h3c];
  assign T650 = T651 == T470;
  assign T651 = idxs[6'h3d];
  assign T2306 = T2307[6'h3d:1'h0];
  assign T2307 = reset ? 64'h0 : T652;
  assign T652 = io_invalidate ? 64'h0 : T653;
  assign T653 = R7 ? T654 : T2308;
  assign T2308 = {2'h0, idxValid};
  assign T654 = T2309 | T655;
  assign T655 = 1'h1 << T42;
  assign T2309 = {2'h0, T656};
  assign T656 = idxValid & T657;
  assign T657 = ~ T658;
  assign T658 = T659;
  assign T659 = {T849, T660};
  assign T660 = {T760, T661};
  assign T661 = {T713, T662};
  assign T662 = {T690, T663};
  assign T663 = {T679, T664};
  assign T664 = {T674, T665};
  assign T665 = T666 != 6'h0;
  assign T666 = pageReplEn & T667;
  assign T667 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T668[3'h5:1'h0];
  assign T668 = 1'h1 << T669;
  assign T669 = tgtPages[6'h0];
  assign T2310 = {T2320, T2311};
  assign T2311 = {T2319, T2312};
  assign T2312 = T2313[1'h1];
  assign T2313 = T2318 | T2314;
  assign T2314 = T2315[1'h1:1'h0];
  assign T2315 = T2317 | T2316;
  assign T2316 = T671[2'h3:1'h0];
  assign T671 = usePageHit ? pageHit : tgtPageRepl;
  assign T2317 = T671[3'h5:3'h4];
  assign T2318 = T2315[2'h3:2'h2];
  assign T2319 = T2318 != 2'h0;
  assign T2320 = T2317 != 2'h0;
  assign T672 = R7 & T673;
  assign T673 = T42 < 6'h3e;
  assign T674 = T675 != 6'h0;
  assign T675 = pageReplEn & T676;
  assign T676 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T677[3'h5:1'h0];
  assign T677 = 1'h1 << T678;
  assign T678 = tgtPages[6'h1];
  assign T679 = {T685, T680};
  assign T680 = T681 != 6'h0;
  assign T681 = pageReplEn & T682;
  assign T682 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T683[3'h5:1'h0];
  assign T683 = 1'h1 << T684;
  assign T684 = tgtPages[6'h2];
  assign T685 = T686 != 6'h0;
  assign T686 = pageReplEn & T687;
  assign T687 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T688[3'h5:1'h0];
  assign T688 = 1'h1 << T689;
  assign T689 = tgtPages[6'h3];
  assign T690 = {T702, T691};
  assign T691 = {T697, T692};
  assign T692 = T693 != 6'h0;
  assign T693 = pageReplEn & T694;
  assign T694 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T695[3'h5:1'h0];
  assign T695 = 1'h1 << T696;
  assign T696 = tgtPages[6'h4];
  assign T697 = T698 != 6'h0;
  assign T698 = pageReplEn & T699;
  assign T699 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T700[3'h5:1'h0];
  assign T700 = 1'h1 << T701;
  assign T701 = tgtPages[6'h5];
  assign T702 = {T708, T703};
  assign T703 = T704 != 6'h0;
  assign T704 = pageReplEn & T705;
  assign T705 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T706[3'h5:1'h0];
  assign T706 = 1'h1 << T707;
  assign T707 = tgtPages[6'h6];
  assign T708 = T709 != 6'h0;
  assign T709 = pageReplEn & T710;
  assign T710 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T711[3'h5:1'h0];
  assign T711 = 1'h1 << T712;
  assign T712 = tgtPages[6'h7];
  assign T713 = {T737, T714};
  assign T714 = {T726, T715};
  assign T715 = {T721, T716};
  assign T716 = T717 != 6'h0;
  assign T717 = pageReplEn & T718;
  assign T718 = idxPagesOH_8 | tgtPagesOH_8;
  assign tgtPagesOH_8 = T719[3'h5:1'h0];
  assign T719 = 1'h1 << T720;
  assign T720 = tgtPages[6'h8];
  assign T721 = T722 != 6'h0;
  assign T722 = pageReplEn & T723;
  assign T723 = idxPagesOH_9 | tgtPagesOH_9;
  assign tgtPagesOH_9 = T724[3'h5:1'h0];
  assign T724 = 1'h1 << T725;
  assign T725 = tgtPages[6'h9];
  assign T726 = {T732, T727};
  assign T727 = T728 != 6'h0;
  assign T728 = pageReplEn & T729;
  assign T729 = idxPagesOH_10 | tgtPagesOH_10;
  assign tgtPagesOH_10 = T730[3'h5:1'h0];
  assign T730 = 1'h1 << T731;
  assign T731 = tgtPages[6'ha];
  assign T732 = T733 != 6'h0;
  assign T733 = pageReplEn & T734;
  assign T734 = idxPagesOH_11 | tgtPagesOH_11;
  assign tgtPagesOH_11 = T735[3'h5:1'h0];
  assign T735 = 1'h1 << T736;
  assign T736 = tgtPages[6'hb];
  assign T737 = {T749, T738};
  assign T738 = {T744, T739};
  assign T739 = T740 != 6'h0;
  assign T740 = pageReplEn & T741;
  assign T741 = idxPagesOH_12 | tgtPagesOH_12;
  assign tgtPagesOH_12 = T742[3'h5:1'h0];
  assign T742 = 1'h1 << T743;
  assign T743 = tgtPages[6'hc];
  assign T744 = T745 != 6'h0;
  assign T745 = pageReplEn & T746;
  assign T746 = idxPagesOH_13 | tgtPagesOH_13;
  assign tgtPagesOH_13 = T747[3'h5:1'h0];
  assign T747 = 1'h1 << T748;
  assign T748 = tgtPages[6'hd];
  assign T749 = {T755, T750};
  assign T750 = T751 != 6'h0;
  assign T751 = pageReplEn & T752;
  assign T752 = idxPagesOH_14 | tgtPagesOH_14;
  assign tgtPagesOH_14 = T753[3'h5:1'h0];
  assign T753 = 1'h1 << T754;
  assign T754 = tgtPages[6'he];
  assign T755 = T756 != 6'h0;
  assign T756 = pageReplEn & T757;
  assign T757 = idxPagesOH_15 | tgtPagesOH_15;
  assign tgtPagesOH_15 = T758[3'h5:1'h0];
  assign T758 = 1'h1 << T759;
  assign T759 = tgtPages[6'hf];
  assign T760 = {T808, T761};
  assign T761 = {T785, T762};
  assign T762 = {T774, T763};
  assign T763 = {T769, T764};
  assign T764 = T765 != 6'h0;
  assign T765 = pageReplEn & T766;
  assign T766 = idxPagesOH_16 | tgtPagesOH_16;
  assign tgtPagesOH_16 = T767[3'h5:1'h0];
  assign T767 = 1'h1 << T768;
  assign T768 = tgtPages[6'h10];
  assign T769 = T770 != 6'h0;
  assign T770 = pageReplEn & T771;
  assign T771 = idxPagesOH_17 | tgtPagesOH_17;
  assign tgtPagesOH_17 = T772[3'h5:1'h0];
  assign T772 = 1'h1 << T773;
  assign T773 = tgtPages[6'h11];
  assign T774 = {T780, T775};
  assign T775 = T776 != 6'h0;
  assign T776 = pageReplEn & T777;
  assign T777 = idxPagesOH_18 | tgtPagesOH_18;
  assign tgtPagesOH_18 = T778[3'h5:1'h0];
  assign T778 = 1'h1 << T779;
  assign T779 = tgtPages[6'h12];
  assign T780 = T781 != 6'h0;
  assign T781 = pageReplEn & T782;
  assign T782 = idxPagesOH_19 | tgtPagesOH_19;
  assign tgtPagesOH_19 = T783[3'h5:1'h0];
  assign T783 = 1'h1 << T784;
  assign T784 = tgtPages[6'h13];
  assign T785 = {T797, T786};
  assign T786 = {T792, T787};
  assign T787 = T788 != 6'h0;
  assign T788 = pageReplEn & T789;
  assign T789 = idxPagesOH_20 | tgtPagesOH_20;
  assign tgtPagesOH_20 = T790[3'h5:1'h0];
  assign T790 = 1'h1 << T791;
  assign T791 = tgtPages[6'h14];
  assign T792 = T793 != 6'h0;
  assign T793 = pageReplEn & T794;
  assign T794 = idxPagesOH_21 | tgtPagesOH_21;
  assign tgtPagesOH_21 = T795[3'h5:1'h0];
  assign T795 = 1'h1 << T796;
  assign T796 = tgtPages[6'h15];
  assign T797 = {T803, T798};
  assign T798 = T799 != 6'h0;
  assign T799 = pageReplEn & T800;
  assign T800 = idxPagesOH_22 | tgtPagesOH_22;
  assign tgtPagesOH_22 = T801[3'h5:1'h0];
  assign T801 = 1'h1 << T802;
  assign T802 = tgtPages[6'h16];
  assign T803 = T804 != 6'h0;
  assign T804 = pageReplEn & T805;
  assign T805 = idxPagesOH_23 | tgtPagesOH_23;
  assign tgtPagesOH_23 = T806[3'h5:1'h0];
  assign T806 = 1'h1 << T807;
  assign T807 = tgtPages[6'h17];
  assign T808 = {T832, T809};
  assign T809 = {T821, T810};
  assign T810 = {T816, T811};
  assign T811 = T812 != 6'h0;
  assign T812 = pageReplEn & T813;
  assign T813 = idxPagesOH_24 | tgtPagesOH_24;
  assign tgtPagesOH_24 = T814[3'h5:1'h0];
  assign T814 = 1'h1 << T815;
  assign T815 = tgtPages[6'h18];
  assign T816 = T817 != 6'h0;
  assign T817 = pageReplEn & T818;
  assign T818 = idxPagesOH_25 | tgtPagesOH_25;
  assign tgtPagesOH_25 = T819[3'h5:1'h0];
  assign T819 = 1'h1 << T820;
  assign T820 = tgtPages[6'h19];
  assign T821 = {T827, T822};
  assign T822 = T823 != 6'h0;
  assign T823 = pageReplEn & T824;
  assign T824 = idxPagesOH_26 | tgtPagesOH_26;
  assign tgtPagesOH_26 = T825[3'h5:1'h0];
  assign T825 = 1'h1 << T826;
  assign T826 = tgtPages[6'h1a];
  assign T827 = T828 != 6'h0;
  assign T828 = pageReplEn & T829;
  assign T829 = idxPagesOH_27 | tgtPagesOH_27;
  assign tgtPagesOH_27 = T830[3'h5:1'h0];
  assign T830 = 1'h1 << T831;
  assign T831 = tgtPages[6'h1b];
  assign T832 = {T844, T833};
  assign T833 = {T839, T834};
  assign T834 = T835 != 6'h0;
  assign T835 = pageReplEn & T836;
  assign T836 = idxPagesOH_28 | tgtPagesOH_28;
  assign tgtPagesOH_28 = T837[3'h5:1'h0];
  assign T837 = 1'h1 << T838;
  assign T838 = tgtPages[6'h1c];
  assign T839 = T840 != 6'h0;
  assign T840 = pageReplEn & T841;
  assign T841 = idxPagesOH_29 | tgtPagesOH_29;
  assign tgtPagesOH_29 = T842[3'h5:1'h0];
  assign T842 = 1'h1 << T843;
  assign T843 = tgtPages[6'h1d];
  assign T844 = T845 != 6'h0;
  assign T845 = pageReplEn & T846;
  assign T846 = idxPagesOH_30 | tgtPagesOH_30;
  assign tgtPagesOH_30 = T847[3'h5:1'h0];
  assign T847 = 1'h1 << T848;
  assign T848 = tgtPages[6'h1e];
  assign T849 = {T945, T850};
  assign T850 = {T898, T851};
  assign T851 = {T875, T852};
  assign T852 = {T864, T853};
  assign T853 = {T859, T854};
  assign T854 = T855 != 6'h0;
  assign T855 = pageReplEn & T856;
  assign T856 = idxPagesOH_31 | tgtPagesOH_31;
  assign tgtPagesOH_31 = T857[3'h5:1'h0];
  assign T857 = 1'h1 << T858;
  assign T858 = tgtPages[6'h1f];
  assign T859 = T860 != 6'h0;
  assign T860 = pageReplEn & T861;
  assign T861 = idxPagesOH_32 | tgtPagesOH_32;
  assign tgtPagesOH_32 = T862[3'h5:1'h0];
  assign T862 = 1'h1 << T863;
  assign T863 = tgtPages[6'h20];
  assign T864 = {T870, T865};
  assign T865 = T866 != 6'h0;
  assign T866 = pageReplEn & T867;
  assign T867 = idxPagesOH_33 | tgtPagesOH_33;
  assign tgtPagesOH_33 = T868[3'h5:1'h0];
  assign T868 = 1'h1 << T869;
  assign T869 = tgtPages[6'h21];
  assign T870 = T871 != 6'h0;
  assign T871 = pageReplEn & T872;
  assign T872 = idxPagesOH_34 | tgtPagesOH_34;
  assign tgtPagesOH_34 = T873[3'h5:1'h0];
  assign T873 = 1'h1 << T874;
  assign T874 = tgtPages[6'h22];
  assign T875 = {T887, T876};
  assign T876 = {T882, T877};
  assign T877 = T878 != 6'h0;
  assign T878 = pageReplEn & T879;
  assign T879 = idxPagesOH_35 | tgtPagesOH_35;
  assign tgtPagesOH_35 = T880[3'h5:1'h0];
  assign T880 = 1'h1 << T881;
  assign T881 = tgtPages[6'h23];
  assign T882 = T883 != 6'h0;
  assign T883 = pageReplEn & T884;
  assign T884 = idxPagesOH_36 | tgtPagesOH_36;
  assign tgtPagesOH_36 = T885[3'h5:1'h0];
  assign T885 = 1'h1 << T886;
  assign T886 = tgtPages[6'h24];
  assign T887 = {T893, T888};
  assign T888 = T889 != 6'h0;
  assign T889 = pageReplEn & T890;
  assign T890 = idxPagesOH_37 | tgtPagesOH_37;
  assign tgtPagesOH_37 = T891[3'h5:1'h0];
  assign T891 = 1'h1 << T892;
  assign T892 = tgtPages[6'h25];
  assign T893 = T894 != 6'h0;
  assign T894 = pageReplEn & T895;
  assign T895 = idxPagesOH_38 | tgtPagesOH_38;
  assign tgtPagesOH_38 = T896[3'h5:1'h0];
  assign T896 = 1'h1 << T897;
  assign T897 = tgtPages[6'h26];
  assign T898 = {T922, T899};
  assign T899 = {T911, T900};
  assign T900 = {T906, T901};
  assign T901 = T902 != 6'h0;
  assign T902 = pageReplEn & T903;
  assign T903 = idxPagesOH_39 | tgtPagesOH_39;
  assign tgtPagesOH_39 = T904[3'h5:1'h0];
  assign T904 = 1'h1 << T905;
  assign T905 = tgtPages[6'h27];
  assign T906 = T907 != 6'h0;
  assign T907 = pageReplEn & T908;
  assign T908 = idxPagesOH_40 | tgtPagesOH_40;
  assign tgtPagesOH_40 = T909[3'h5:1'h0];
  assign T909 = 1'h1 << T910;
  assign T910 = tgtPages[6'h28];
  assign T911 = {T917, T912};
  assign T912 = T913 != 6'h0;
  assign T913 = pageReplEn & T914;
  assign T914 = idxPagesOH_41 | tgtPagesOH_41;
  assign tgtPagesOH_41 = T915[3'h5:1'h0];
  assign T915 = 1'h1 << T916;
  assign T916 = tgtPages[6'h29];
  assign T917 = T918 != 6'h0;
  assign T918 = pageReplEn & T919;
  assign T919 = idxPagesOH_42 | tgtPagesOH_42;
  assign tgtPagesOH_42 = T920[3'h5:1'h0];
  assign T920 = 1'h1 << T921;
  assign T921 = tgtPages[6'h2a];
  assign T922 = {T934, T923};
  assign T923 = {T929, T924};
  assign T924 = T925 != 6'h0;
  assign T925 = pageReplEn & T926;
  assign T926 = idxPagesOH_43 | tgtPagesOH_43;
  assign tgtPagesOH_43 = T927[3'h5:1'h0];
  assign T927 = 1'h1 << T928;
  assign T928 = tgtPages[6'h2b];
  assign T929 = T930 != 6'h0;
  assign T930 = pageReplEn & T931;
  assign T931 = idxPagesOH_44 | tgtPagesOH_44;
  assign tgtPagesOH_44 = T932[3'h5:1'h0];
  assign T932 = 1'h1 << T933;
  assign T933 = tgtPages[6'h2c];
  assign T934 = {T940, T935};
  assign T935 = T936 != 6'h0;
  assign T936 = pageReplEn & T937;
  assign T937 = idxPagesOH_45 | tgtPagesOH_45;
  assign tgtPagesOH_45 = T938[3'h5:1'h0];
  assign T938 = 1'h1 << T939;
  assign T939 = tgtPages[6'h2d];
  assign T940 = T941 != 6'h0;
  assign T941 = pageReplEn & T942;
  assign T942 = idxPagesOH_46 | tgtPagesOH_46;
  assign tgtPagesOH_46 = T943[3'h5:1'h0];
  assign T943 = 1'h1 << T944;
  assign T944 = tgtPages[6'h2e];
  assign T945 = {T993, T946};
  assign T946 = {T970, T947};
  assign T947 = {T959, T948};
  assign T948 = {T954, T949};
  assign T949 = T950 != 6'h0;
  assign T950 = pageReplEn & T951;
  assign T951 = idxPagesOH_47 | tgtPagesOH_47;
  assign tgtPagesOH_47 = T952[3'h5:1'h0];
  assign T952 = 1'h1 << T953;
  assign T953 = tgtPages[6'h2f];
  assign T954 = T955 != 6'h0;
  assign T955 = pageReplEn & T956;
  assign T956 = idxPagesOH_48 | tgtPagesOH_48;
  assign tgtPagesOH_48 = T957[3'h5:1'h0];
  assign T957 = 1'h1 << T958;
  assign T958 = tgtPages[6'h30];
  assign T959 = {T965, T960};
  assign T960 = T961 != 6'h0;
  assign T961 = pageReplEn & T962;
  assign T962 = idxPagesOH_49 | tgtPagesOH_49;
  assign tgtPagesOH_49 = T963[3'h5:1'h0];
  assign T963 = 1'h1 << T964;
  assign T964 = tgtPages[6'h31];
  assign T965 = T966 != 6'h0;
  assign T966 = pageReplEn & T967;
  assign T967 = idxPagesOH_50 | tgtPagesOH_50;
  assign tgtPagesOH_50 = T968[3'h5:1'h0];
  assign T968 = 1'h1 << T969;
  assign T969 = tgtPages[6'h32];
  assign T970 = {T982, T971};
  assign T971 = {T977, T972};
  assign T972 = T973 != 6'h0;
  assign T973 = pageReplEn & T974;
  assign T974 = idxPagesOH_51 | tgtPagesOH_51;
  assign tgtPagesOH_51 = T975[3'h5:1'h0];
  assign T975 = 1'h1 << T976;
  assign T976 = tgtPages[6'h33];
  assign T977 = T978 != 6'h0;
  assign T978 = pageReplEn & T979;
  assign T979 = idxPagesOH_52 | tgtPagesOH_52;
  assign tgtPagesOH_52 = T980[3'h5:1'h0];
  assign T980 = 1'h1 << T981;
  assign T981 = tgtPages[6'h34];
  assign T982 = {T988, T983};
  assign T983 = T984 != 6'h0;
  assign T984 = pageReplEn & T985;
  assign T985 = idxPagesOH_53 | tgtPagesOH_53;
  assign tgtPagesOH_53 = T986[3'h5:1'h0];
  assign T986 = 1'h1 << T987;
  assign T987 = tgtPages[6'h35];
  assign T988 = T989 != 6'h0;
  assign T989 = pageReplEn & T990;
  assign T990 = idxPagesOH_54 | tgtPagesOH_54;
  assign tgtPagesOH_54 = T991[3'h5:1'h0];
  assign T991 = 1'h1 << T992;
  assign T992 = tgtPages[6'h36];
  assign T993 = {T1017, T994};
  assign T994 = {T1006, T995};
  assign T995 = {T1001, T996};
  assign T996 = T997 != 6'h0;
  assign T997 = pageReplEn & T998;
  assign T998 = idxPagesOH_55 | tgtPagesOH_55;
  assign tgtPagesOH_55 = T999[3'h5:1'h0];
  assign T999 = 1'h1 << T1000;
  assign T1000 = tgtPages[6'h37];
  assign T1001 = T1002 != 6'h0;
  assign T1002 = pageReplEn & T1003;
  assign T1003 = idxPagesOH_56 | tgtPagesOH_56;
  assign tgtPagesOH_56 = T1004[3'h5:1'h0];
  assign T1004 = 1'h1 << T1005;
  assign T1005 = tgtPages[6'h38];
  assign T1006 = {T1012, T1007};
  assign T1007 = T1008 != 6'h0;
  assign T1008 = pageReplEn & T1009;
  assign T1009 = idxPagesOH_57 | tgtPagesOH_57;
  assign tgtPagesOH_57 = T1010[3'h5:1'h0];
  assign T1010 = 1'h1 << T1011;
  assign T1011 = tgtPages[6'h39];
  assign T1012 = T1013 != 6'h0;
  assign T1013 = pageReplEn & T1014;
  assign T1014 = idxPagesOH_58 | tgtPagesOH_58;
  assign tgtPagesOH_58 = T1015[3'h5:1'h0];
  assign T1015 = 1'h1 << T1016;
  assign T1016 = tgtPages[6'h3a];
  assign T1017 = {T1029, T1018};
  assign T1018 = {T1024, T1019};
  assign T1019 = T1020 != 6'h0;
  assign T1020 = pageReplEn & T1021;
  assign T1021 = idxPagesOH_59 | tgtPagesOH_59;
  assign tgtPagesOH_59 = T1022[3'h5:1'h0];
  assign T1022 = 1'h1 << T1023;
  assign T1023 = tgtPages[6'h3b];
  assign T1024 = T1025 != 6'h0;
  assign T1025 = pageReplEn & T1026;
  assign T1026 = idxPagesOH_60 | tgtPagesOH_60;
  assign tgtPagesOH_60 = T1027[3'h5:1'h0];
  assign T1027 = 1'h1 << T1028;
  assign T1028 = tgtPages[6'h3c];
  assign T1029 = T1030 != 6'h0;
  assign T1030 = pageReplEn & T1031;
  assign T1031 = idxPagesOH_61 | tgtPagesOH_61;
  assign tgtPagesOH_61 = T1032[3'h5:1'h0];
  assign T1032 = 1'h1 << T1033;
  assign T1033 = tgtPages[6'h3d];
  assign T1034 = T1040 | T1035;
  assign T1035 = T1039 ? isJump_60 : 1'h0;
  assign T1036 = T1037 ? R36 : isJump_60;
  assign T1037 = R7 & T1038;
  assign T1038 = T40[6'h3c];
  assign T1039 = hits[6'h3c];
  assign T1040 = T1046 | T1041;
  assign T1041 = T1045 ? isJump_59 : 1'h0;
  assign T1042 = T1043 ? R36 : isJump_59;
  assign T1043 = R7 & T1044;
  assign T1044 = T40[6'h3b];
  assign T1045 = hits[6'h3b];
  assign T1046 = T1052 | T1047;
  assign T1047 = T1051 ? isJump_58 : 1'h0;
  assign T1048 = T1049 ? R36 : isJump_58;
  assign T1049 = R7 & T1050;
  assign T1050 = T40[6'h3a];
  assign T1051 = hits[6'h3a];
  assign T1052 = T1058 | T1053;
  assign T1053 = T1057 ? isJump_57 : 1'h0;
  assign T1054 = T1055 ? R36 : isJump_57;
  assign T1055 = R7 & T1056;
  assign T1056 = T40[6'h39];
  assign T1057 = hits[6'h39];
  assign T1058 = T1064 | T1059;
  assign T1059 = T1063 ? isJump_56 : 1'h0;
  assign T1060 = T1061 ? R36 : isJump_56;
  assign T1061 = R7 & T1062;
  assign T1062 = T40[6'h38];
  assign T1063 = hits[6'h38];
  assign T1064 = T1070 | T1065;
  assign T1065 = T1069 ? isJump_55 : 1'h0;
  assign T1066 = T1067 ? R36 : isJump_55;
  assign T1067 = R7 & T1068;
  assign T1068 = T40[6'h37];
  assign T1069 = hits[6'h37];
  assign T1070 = T1076 | T1071;
  assign T1071 = T1075 ? isJump_54 : 1'h0;
  assign T1072 = T1073 ? R36 : isJump_54;
  assign T1073 = R7 & T1074;
  assign T1074 = T40[6'h36];
  assign T1075 = hits[6'h36];
  assign T1076 = T1082 | T1077;
  assign T1077 = T1081 ? isJump_53 : 1'h0;
  assign T1078 = T1079 ? R36 : isJump_53;
  assign T1079 = R7 & T1080;
  assign T1080 = T40[6'h35];
  assign T1081 = hits[6'h35];
  assign T1082 = T1088 | T1083;
  assign T1083 = T1087 ? isJump_52 : 1'h0;
  assign T1084 = T1085 ? R36 : isJump_52;
  assign T1085 = R7 & T1086;
  assign T1086 = T40[6'h34];
  assign T1087 = hits[6'h34];
  assign T1088 = T1094 | T1089;
  assign T1089 = T1093 ? isJump_51 : 1'h0;
  assign T1090 = T1091 ? R36 : isJump_51;
  assign T1091 = R7 & T1092;
  assign T1092 = T40[6'h33];
  assign T1093 = hits[6'h33];
  assign T1094 = T1100 | T1095;
  assign T1095 = T1099 ? isJump_50 : 1'h0;
  assign T1096 = T1097 ? R36 : isJump_50;
  assign T1097 = R7 & T1098;
  assign T1098 = T40[6'h32];
  assign T1099 = hits[6'h32];
  assign T1100 = T1106 | T1101;
  assign T1101 = T1105 ? isJump_49 : 1'h0;
  assign T1102 = T1103 ? R36 : isJump_49;
  assign T1103 = R7 & T1104;
  assign T1104 = T40[6'h31];
  assign T1105 = hits[6'h31];
  assign T1106 = T1112 | T1107;
  assign T1107 = T1111 ? isJump_48 : 1'h0;
  assign T1108 = T1109 ? R36 : isJump_48;
  assign T1109 = R7 & T1110;
  assign T1110 = T40[6'h30];
  assign T1111 = hits[6'h30];
  assign T1112 = T1118 | T1113;
  assign T1113 = T1117 ? isJump_47 : 1'h0;
  assign T1114 = T1115 ? R36 : isJump_47;
  assign T1115 = R7 & T1116;
  assign T1116 = T40[6'h2f];
  assign T1117 = hits[6'h2f];
  assign T1118 = T1124 | T1119;
  assign T1119 = T1123 ? isJump_46 : 1'h0;
  assign T1120 = T1121 ? R36 : isJump_46;
  assign T1121 = R7 & T1122;
  assign T1122 = T40[6'h2e];
  assign T1123 = hits[6'h2e];
  assign T1124 = T1130 | T1125;
  assign T1125 = T1129 ? isJump_45 : 1'h0;
  assign T1126 = T1127 ? R36 : isJump_45;
  assign T1127 = R7 & T1128;
  assign T1128 = T40[6'h2d];
  assign T1129 = hits[6'h2d];
  assign T1130 = T1136 | T1131;
  assign T1131 = T1135 ? isJump_44 : 1'h0;
  assign T1132 = T1133 ? R36 : isJump_44;
  assign T1133 = R7 & T1134;
  assign T1134 = T40[6'h2c];
  assign T1135 = hits[6'h2c];
  assign T1136 = T1142 | T1137;
  assign T1137 = T1141 ? isJump_43 : 1'h0;
  assign T1138 = T1139 ? R36 : isJump_43;
  assign T1139 = R7 & T1140;
  assign T1140 = T40[6'h2b];
  assign T1141 = hits[6'h2b];
  assign T1142 = T1148 | T1143;
  assign T1143 = T1147 ? isJump_42 : 1'h0;
  assign T1144 = T1145 ? R36 : isJump_42;
  assign T1145 = R7 & T1146;
  assign T1146 = T40[6'h2a];
  assign T1147 = hits[6'h2a];
  assign T1148 = T1154 | T1149;
  assign T1149 = T1153 ? isJump_41 : 1'h0;
  assign T1150 = T1151 ? R36 : isJump_41;
  assign T1151 = R7 & T1152;
  assign T1152 = T40[6'h29];
  assign T1153 = hits[6'h29];
  assign T1154 = T1160 | T1155;
  assign T1155 = T1159 ? isJump_40 : 1'h0;
  assign T1156 = T1157 ? R36 : isJump_40;
  assign T1157 = R7 & T1158;
  assign T1158 = T40[6'h28];
  assign T1159 = hits[6'h28];
  assign T1160 = T1166 | T1161;
  assign T1161 = T1165 ? isJump_39 : 1'h0;
  assign T1162 = T1163 ? R36 : isJump_39;
  assign T1163 = R7 & T1164;
  assign T1164 = T40[6'h27];
  assign T1165 = hits[6'h27];
  assign T1166 = T1172 | T1167;
  assign T1167 = T1171 ? isJump_38 : 1'h0;
  assign T1168 = T1169 ? R36 : isJump_38;
  assign T1169 = R7 & T1170;
  assign T1170 = T40[6'h26];
  assign T1171 = hits[6'h26];
  assign T1172 = T1178 | T1173;
  assign T1173 = T1177 ? isJump_37 : 1'h0;
  assign T1174 = T1175 ? R36 : isJump_37;
  assign T1175 = R7 & T1176;
  assign T1176 = T40[6'h25];
  assign T1177 = hits[6'h25];
  assign T1178 = T1184 | T1179;
  assign T1179 = T1183 ? isJump_36 : 1'h0;
  assign T1180 = T1181 ? R36 : isJump_36;
  assign T1181 = R7 & T1182;
  assign T1182 = T40[6'h24];
  assign T1183 = hits[6'h24];
  assign T1184 = T1190 | T1185;
  assign T1185 = T1189 ? isJump_35 : 1'h0;
  assign T1186 = T1187 ? R36 : isJump_35;
  assign T1187 = R7 & T1188;
  assign T1188 = T40[6'h23];
  assign T1189 = hits[6'h23];
  assign T1190 = T1196 | T1191;
  assign T1191 = T1195 ? isJump_34 : 1'h0;
  assign T1192 = T1193 ? R36 : isJump_34;
  assign T1193 = R7 & T1194;
  assign T1194 = T40[6'h22];
  assign T1195 = hits[6'h22];
  assign T1196 = T1202 | T1197;
  assign T1197 = T1201 ? isJump_33 : 1'h0;
  assign T1198 = T1199 ? R36 : isJump_33;
  assign T1199 = R7 & T1200;
  assign T1200 = T40[6'h21];
  assign T1201 = hits[6'h21];
  assign T1202 = T1208 | T1203;
  assign T1203 = T1207 ? isJump_32 : 1'h0;
  assign T1204 = T1205 ? R36 : isJump_32;
  assign T1205 = R7 & T1206;
  assign T1206 = T40[6'h20];
  assign T1207 = hits[6'h20];
  assign T1208 = T1214 | T1209;
  assign T1209 = T1213 ? isJump_31 : 1'h0;
  assign T1210 = T1211 ? R36 : isJump_31;
  assign T1211 = R7 & T1212;
  assign T1212 = T40[5'h1f];
  assign T1213 = hits[5'h1f];
  assign T1214 = T1220 | T1215;
  assign T1215 = T1219 ? isJump_30 : 1'h0;
  assign T1216 = T1217 ? R36 : isJump_30;
  assign T1217 = R7 & T1218;
  assign T1218 = T40[5'h1e];
  assign T1219 = hits[5'h1e];
  assign T1220 = T1226 | T1221;
  assign T1221 = T1225 ? isJump_29 : 1'h0;
  assign T1222 = T1223 ? R36 : isJump_29;
  assign T1223 = R7 & T1224;
  assign T1224 = T40[5'h1d];
  assign T1225 = hits[5'h1d];
  assign T1226 = T1232 | T1227;
  assign T1227 = T1231 ? isJump_28 : 1'h0;
  assign T1228 = T1229 ? R36 : isJump_28;
  assign T1229 = R7 & T1230;
  assign T1230 = T40[5'h1c];
  assign T1231 = hits[5'h1c];
  assign T1232 = T1238 | T1233;
  assign T1233 = T1237 ? isJump_27 : 1'h0;
  assign T1234 = T1235 ? R36 : isJump_27;
  assign T1235 = R7 & T1236;
  assign T1236 = T40[5'h1b];
  assign T1237 = hits[5'h1b];
  assign T1238 = T1244 | T1239;
  assign T1239 = T1243 ? isJump_26 : 1'h0;
  assign T1240 = T1241 ? R36 : isJump_26;
  assign T1241 = R7 & T1242;
  assign T1242 = T40[5'h1a];
  assign T1243 = hits[5'h1a];
  assign T1244 = T1250 | T1245;
  assign T1245 = T1249 ? isJump_25 : 1'h0;
  assign T1246 = T1247 ? R36 : isJump_25;
  assign T1247 = R7 & T1248;
  assign T1248 = T40[5'h19];
  assign T1249 = hits[5'h19];
  assign T1250 = T1256 | T1251;
  assign T1251 = T1255 ? isJump_24 : 1'h0;
  assign T1252 = T1253 ? R36 : isJump_24;
  assign T1253 = R7 & T1254;
  assign T1254 = T40[5'h18];
  assign T1255 = hits[5'h18];
  assign T1256 = T1262 | T1257;
  assign T1257 = T1261 ? isJump_23 : 1'h0;
  assign T1258 = T1259 ? R36 : isJump_23;
  assign T1259 = R7 & T1260;
  assign T1260 = T40[5'h17];
  assign T1261 = hits[5'h17];
  assign T1262 = T1268 | T1263;
  assign T1263 = T1267 ? isJump_22 : 1'h0;
  assign T1264 = T1265 ? R36 : isJump_22;
  assign T1265 = R7 & T1266;
  assign T1266 = T40[5'h16];
  assign T1267 = hits[5'h16];
  assign T1268 = T1274 | T1269;
  assign T1269 = T1273 ? isJump_21 : 1'h0;
  assign T1270 = T1271 ? R36 : isJump_21;
  assign T1271 = R7 & T1272;
  assign T1272 = T40[5'h15];
  assign T1273 = hits[5'h15];
  assign T1274 = T1280 | T1275;
  assign T1275 = T1279 ? isJump_20 : 1'h0;
  assign T1276 = T1277 ? R36 : isJump_20;
  assign T1277 = R7 & T1278;
  assign T1278 = T40[5'h14];
  assign T1279 = hits[5'h14];
  assign T1280 = T1286 | T1281;
  assign T1281 = T1285 ? isJump_19 : 1'h0;
  assign T1282 = T1283 ? R36 : isJump_19;
  assign T1283 = R7 & T1284;
  assign T1284 = T40[5'h13];
  assign T1285 = hits[5'h13];
  assign T1286 = T1292 | T1287;
  assign T1287 = T1291 ? isJump_18 : 1'h0;
  assign T1288 = T1289 ? R36 : isJump_18;
  assign T1289 = R7 & T1290;
  assign T1290 = T40[5'h12];
  assign T1291 = hits[5'h12];
  assign T1292 = T1298 | T1293;
  assign T1293 = T1297 ? isJump_17 : 1'h0;
  assign T1294 = T1295 ? R36 : isJump_17;
  assign T1295 = R7 & T1296;
  assign T1296 = T40[5'h11];
  assign T1297 = hits[5'h11];
  assign T1298 = T1304 | T1299;
  assign T1299 = T1303 ? isJump_16 : 1'h0;
  assign T1300 = T1301 ? R36 : isJump_16;
  assign T1301 = R7 & T1302;
  assign T1302 = T40[5'h10];
  assign T1303 = hits[5'h10];
  assign T1304 = T1310 | T1305;
  assign T1305 = T1309 ? isJump_15 : 1'h0;
  assign T1306 = T1307 ? R36 : isJump_15;
  assign T1307 = R7 & T1308;
  assign T1308 = T40[4'hf];
  assign T1309 = hits[4'hf];
  assign T1310 = T1316 | T1311;
  assign T1311 = T1315 ? isJump_14 : 1'h0;
  assign T1312 = T1313 ? R36 : isJump_14;
  assign T1313 = R7 & T1314;
  assign T1314 = T40[4'he];
  assign T1315 = hits[4'he];
  assign T1316 = T1322 | T1317;
  assign T1317 = T1321 ? isJump_13 : 1'h0;
  assign T1318 = T1319 ? R36 : isJump_13;
  assign T1319 = R7 & T1320;
  assign T1320 = T40[4'hd];
  assign T1321 = hits[4'hd];
  assign T1322 = T1328 | T1323;
  assign T1323 = T1327 ? isJump_12 : 1'h0;
  assign T1324 = T1325 ? R36 : isJump_12;
  assign T1325 = R7 & T1326;
  assign T1326 = T40[4'hc];
  assign T1327 = hits[4'hc];
  assign T1328 = T1334 | T1329;
  assign T1329 = T1333 ? isJump_11 : 1'h0;
  assign T1330 = T1331 ? R36 : isJump_11;
  assign T1331 = R7 & T1332;
  assign T1332 = T40[4'hb];
  assign T1333 = hits[4'hb];
  assign T1334 = T1340 | T1335;
  assign T1335 = T1339 ? isJump_10 : 1'h0;
  assign T1336 = T1337 ? R36 : isJump_10;
  assign T1337 = R7 & T1338;
  assign T1338 = T40[4'ha];
  assign T1339 = hits[4'ha];
  assign T1340 = T1346 | T1341;
  assign T1341 = T1345 ? isJump_9 : 1'h0;
  assign T1342 = T1343 ? R36 : isJump_9;
  assign T1343 = R7 & T1344;
  assign T1344 = T40[4'h9];
  assign T1345 = hits[4'h9];
  assign T1346 = T1352 | T1347;
  assign T1347 = T1351 ? isJump_8 : 1'h0;
  assign T1348 = T1349 ? R36 : isJump_8;
  assign T1349 = R7 & T1350;
  assign T1350 = T40[4'h8];
  assign T1351 = hits[4'h8];
  assign T1352 = T1358 | T1353;
  assign T1353 = T1357 ? isJump_7 : 1'h0;
  assign T1354 = T1355 ? R36 : isJump_7;
  assign T1355 = R7 & T1356;
  assign T1356 = T40[3'h7];
  assign T1357 = hits[3'h7];
  assign T1358 = T1364 | T1359;
  assign T1359 = T1363 ? isJump_6 : 1'h0;
  assign T1360 = T1361 ? R36 : isJump_6;
  assign T1361 = R7 & T1362;
  assign T1362 = T40[3'h6];
  assign T1363 = hits[3'h6];
  assign T1364 = T1370 | T1365;
  assign T1365 = T1369 ? isJump_5 : 1'h0;
  assign T1366 = T1367 ? R36 : isJump_5;
  assign T1367 = R7 & T1368;
  assign T1368 = T40[3'h5];
  assign T1369 = hits[3'h5];
  assign T1370 = T1376 | T1371;
  assign T1371 = T1375 ? isJump_4 : 1'h0;
  assign T1372 = T1373 ? R36 : isJump_4;
  assign T1373 = R7 & T1374;
  assign T1374 = T40[3'h4];
  assign T1375 = hits[3'h4];
  assign T1376 = T1382 | T1377;
  assign T1377 = T1381 ? isJump_3 : 1'h0;
  assign T1378 = T1379 ? R36 : isJump_3;
  assign T1379 = R7 & T1380;
  assign T1380 = T40[2'h3];
  assign T1381 = hits[2'h3];
  assign T1382 = T1388 | T1383;
  assign T1383 = T1387 ? isJump_2 : 1'h0;
  assign T1384 = T1385 ? R36 : isJump_2;
  assign T1385 = R7 & T1386;
  assign T1386 = T40[2'h2];
  assign T1387 = hits[2'h2];
  assign T1388 = T1394 | T1389;
  assign T1389 = T1393 ? isJump_1 : 1'h0;
  assign T1390 = T1391 ? R36 : isJump_1;
  assign T1391 = R7 & T1392;
  assign T1392 = T40[1'h1];
  assign T1393 = hits[1'h1];
  assign T1394 = T1398 ? isJump_0 : 1'h0;
  assign T1395 = T1396 ? R36 : isJump_0;
  assign T1396 = R7 & T1397;
  assign T1397 = T40[1'h0];
  assign T1398 = hits[1'h0];
  assign T1399 = io_req_valid & io_resp_valid;
  assign T1400 = {io_bht_update_bits_taken, T1401};
  assign T1401 = io_bht_update_bits_prediction_bits_bht_history[3'h6:1'h1];
  assign T1402 = T21 & io_bht_update_bits_mispredict;
  assign T1403 = io_req_bits_addr[4'h8:2'h2];
  assign io_resp_bits_bht_history = T1404;
  assign T1404 = R25;
  assign io_resp_bits_entry = T2321;
  assign T2321 = {T2346, T2322};
  assign T2322 = {T2345, T2323};
  assign T2323 = {T2344, T2324};
  assign T2324 = {T2343, T2325};
  assign T2325 = {T2342, T2326};
  assign T2326 = T2327[1'h1];
  assign T2327 = T2341 | T2328;
  assign T2328 = T2329[1'h1:1'h0];
  assign T2329 = T2340 | T2330;
  assign T2330 = T2331[2'h3:1'h0];
  assign T2331 = T2339 | T2332;
  assign T2332 = T2333[3'h7:1'h0];
  assign T2333 = T2338 | T2334;
  assign T2334 = T2335[4'hf:1'h0];
  assign T2335 = T2337 | T2336;
  assign T2336 = hits[5'h1f:1'h0];
  assign T2337 = hits[6'h3d:6'h20];
  assign T2338 = T2335[5'h1f:5'h10];
  assign T2339 = T2333[4'hf:4'h8];
  assign T2340 = T2331[3'h7:3'h4];
  assign T2341 = T2329[2'h3:2'h2];
  assign T2342 = T2341 != 2'h0;
  assign T2343 = T2340 != 4'h0;
  assign T2344 = T2339 != 8'h0;
  assign T2345 = T2338 != 16'h0;
  assign T2346 = T2337 != 30'h0;
  assign io_resp_bits_target = T1406;
  assign T1406 = T2278 ? io_ras_update_bits_returnAddr : T1407;
  assign T1407 = T1900 ? T1867 : T1408;
  assign T1408 = {T1659, T1409};
  assign T1409 = T1416 | T1410;
  assign T1410 = T1415 ? T1411 : 12'h0;
  assign T1411 = tgts[6'h3d];
  assign T2347 = io_req_bits_addr[4'hb:1'h0];
  assign T1413 = R7 & T1414;
  assign T1414 = T42 < 6'h3e;
  assign T1415 = hits[6'h3d];
  assign T1416 = T1420 | T1417;
  assign T1417 = T1419 ? T1418 : 12'h0;
  assign T1418 = tgts[6'h3c];
  assign T1419 = hits[6'h3c];
  assign T1420 = T1424 | T1421;
  assign T1421 = T1423 ? T1422 : 12'h0;
  assign T1422 = tgts[6'h3b];
  assign T1423 = hits[6'h3b];
  assign T1424 = T1428 | T1425;
  assign T1425 = T1427 ? T1426 : 12'h0;
  assign T1426 = tgts[6'h3a];
  assign T1427 = hits[6'h3a];
  assign T1428 = T1432 | T1429;
  assign T1429 = T1431 ? T1430 : 12'h0;
  assign T1430 = tgts[6'h39];
  assign T1431 = hits[6'h39];
  assign T1432 = T1436 | T1433;
  assign T1433 = T1435 ? T1434 : 12'h0;
  assign T1434 = tgts[6'h38];
  assign T1435 = hits[6'h38];
  assign T1436 = T1440 | T1437;
  assign T1437 = T1439 ? T1438 : 12'h0;
  assign T1438 = tgts[6'h37];
  assign T1439 = hits[6'h37];
  assign T1440 = T1444 | T1441;
  assign T1441 = T1443 ? T1442 : 12'h0;
  assign T1442 = tgts[6'h36];
  assign T1443 = hits[6'h36];
  assign T1444 = T1448 | T1445;
  assign T1445 = T1447 ? T1446 : 12'h0;
  assign T1446 = tgts[6'h35];
  assign T1447 = hits[6'h35];
  assign T1448 = T1452 | T1449;
  assign T1449 = T1451 ? T1450 : 12'h0;
  assign T1450 = tgts[6'h34];
  assign T1451 = hits[6'h34];
  assign T1452 = T1456 | T1453;
  assign T1453 = T1455 ? T1454 : 12'h0;
  assign T1454 = tgts[6'h33];
  assign T1455 = hits[6'h33];
  assign T1456 = T1460 | T1457;
  assign T1457 = T1459 ? T1458 : 12'h0;
  assign T1458 = tgts[6'h32];
  assign T1459 = hits[6'h32];
  assign T1460 = T1464 | T1461;
  assign T1461 = T1463 ? T1462 : 12'h0;
  assign T1462 = tgts[6'h31];
  assign T1463 = hits[6'h31];
  assign T1464 = T1468 | T1465;
  assign T1465 = T1467 ? T1466 : 12'h0;
  assign T1466 = tgts[6'h30];
  assign T1467 = hits[6'h30];
  assign T1468 = T1472 | T1469;
  assign T1469 = T1471 ? T1470 : 12'h0;
  assign T1470 = tgts[6'h2f];
  assign T1471 = hits[6'h2f];
  assign T1472 = T1476 | T1473;
  assign T1473 = T1475 ? T1474 : 12'h0;
  assign T1474 = tgts[6'h2e];
  assign T1475 = hits[6'h2e];
  assign T1476 = T1480 | T1477;
  assign T1477 = T1479 ? T1478 : 12'h0;
  assign T1478 = tgts[6'h2d];
  assign T1479 = hits[6'h2d];
  assign T1480 = T1484 | T1481;
  assign T1481 = T1483 ? T1482 : 12'h0;
  assign T1482 = tgts[6'h2c];
  assign T1483 = hits[6'h2c];
  assign T1484 = T1488 | T1485;
  assign T1485 = T1487 ? T1486 : 12'h0;
  assign T1486 = tgts[6'h2b];
  assign T1487 = hits[6'h2b];
  assign T1488 = T1492 | T1489;
  assign T1489 = T1491 ? T1490 : 12'h0;
  assign T1490 = tgts[6'h2a];
  assign T1491 = hits[6'h2a];
  assign T1492 = T1496 | T1493;
  assign T1493 = T1495 ? T1494 : 12'h0;
  assign T1494 = tgts[6'h29];
  assign T1495 = hits[6'h29];
  assign T1496 = T1500 | T1497;
  assign T1497 = T1499 ? T1498 : 12'h0;
  assign T1498 = tgts[6'h28];
  assign T1499 = hits[6'h28];
  assign T1500 = T1504 | T1501;
  assign T1501 = T1503 ? T1502 : 12'h0;
  assign T1502 = tgts[6'h27];
  assign T1503 = hits[6'h27];
  assign T1504 = T1508 | T1505;
  assign T1505 = T1507 ? T1506 : 12'h0;
  assign T1506 = tgts[6'h26];
  assign T1507 = hits[6'h26];
  assign T1508 = T1512 | T1509;
  assign T1509 = T1511 ? T1510 : 12'h0;
  assign T1510 = tgts[6'h25];
  assign T1511 = hits[6'h25];
  assign T1512 = T1516 | T1513;
  assign T1513 = T1515 ? T1514 : 12'h0;
  assign T1514 = tgts[6'h24];
  assign T1515 = hits[6'h24];
  assign T1516 = T1520 | T1517;
  assign T1517 = T1519 ? T1518 : 12'h0;
  assign T1518 = tgts[6'h23];
  assign T1519 = hits[6'h23];
  assign T1520 = T1524 | T1521;
  assign T1521 = T1523 ? T1522 : 12'h0;
  assign T1522 = tgts[6'h22];
  assign T1523 = hits[6'h22];
  assign T1524 = T1528 | T1525;
  assign T1525 = T1527 ? T1526 : 12'h0;
  assign T1526 = tgts[6'h21];
  assign T1527 = hits[6'h21];
  assign T1528 = T1532 | T1529;
  assign T1529 = T1531 ? T1530 : 12'h0;
  assign T1530 = tgts[6'h20];
  assign T1531 = hits[6'h20];
  assign T1532 = T1536 | T1533;
  assign T1533 = T1535 ? T1534 : 12'h0;
  assign T1534 = tgts[6'h1f];
  assign T1535 = hits[5'h1f];
  assign T1536 = T1540 | T1537;
  assign T1537 = T1539 ? T1538 : 12'h0;
  assign T1538 = tgts[6'h1e];
  assign T1539 = hits[5'h1e];
  assign T1540 = T1544 | T1541;
  assign T1541 = T1543 ? T1542 : 12'h0;
  assign T1542 = tgts[6'h1d];
  assign T1543 = hits[5'h1d];
  assign T1544 = T1548 | T1545;
  assign T1545 = T1547 ? T1546 : 12'h0;
  assign T1546 = tgts[6'h1c];
  assign T1547 = hits[5'h1c];
  assign T1548 = T1552 | T1549;
  assign T1549 = T1551 ? T1550 : 12'h0;
  assign T1550 = tgts[6'h1b];
  assign T1551 = hits[5'h1b];
  assign T1552 = T1556 | T1553;
  assign T1553 = T1555 ? T1554 : 12'h0;
  assign T1554 = tgts[6'h1a];
  assign T1555 = hits[5'h1a];
  assign T1556 = T1560 | T1557;
  assign T1557 = T1559 ? T1558 : 12'h0;
  assign T1558 = tgts[6'h19];
  assign T1559 = hits[5'h19];
  assign T1560 = T1564 | T1561;
  assign T1561 = T1563 ? T1562 : 12'h0;
  assign T1562 = tgts[6'h18];
  assign T1563 = hits[5'h18];
  assign T1564 = T1568 | T1565;
  assign T1565 = T1567 ? T1566 : 12'h0;
  assign T1566 = tgts[6'h17];
  assign T1567 = hits[5'h17];
  assign T1568 = T1572 | T1569;
  assign T1569 = T1571 ? T1570 : 12'h0;
  assign T1570 = tgts[6'h16];
  assign T1571 = hits[5'h16];
  assign T1572 = T1576 | T1573;
  assign T1573 = T1575 ? T1574 : 12'h0;
  assign T1574 = tgts[6'h15];
  assign T1575 = hits[5'h15];
  assign T1576 = T1580 | T1577;
  assign T1577 = T1579 ? T1578 : 12'h0;
  assign T1578 = tgts[6'h14];
  assign T1579 = hits[5'h14];
  assign T1580 = T1584 | T1581;
  assign T1581 = T1583 ? T1582 : 12'h0;
  assign T1582 = tgts[6'h13];
  assign T1583 = hits[5'h13];
  assign T1584 = T1588 | T1585;
  assign T1585 = T1587 ? T1586 : 12'h0;
  assign T1586 = tgts[6'h12];
  assign T1587 = hits[5'h12];
  assign T1588 = T1592 | T1589;
  assign T1589 = T1591 ? T1590 : 12'h0;
  assign T1590 = tgts[6'h11];
  assign T1591 = hits[5'h11];
  assign T1592 = T1596 | T1593;
  assign T1593 = T1595 ? T1594 : 12'h0;
  assign T1594 = tgts[6'h10];
  assign T1595 = hits[5'h10];
  assign T1596 = T1600 | T1597;
  assign T1597 = T1599 ? T1598 : 12'h0;
  assign T1598 = tgts[6'hf];
  assign T1599 = hits[4'hf];
  assign T1600 = T1604 | T1601;
  assign T1601 = T1603 ? T1602 : 12'h0;
  assign T1602 = tgts[6'he];
  assign T1603 = hits[4'he];
  assign T1604 = T1608 | T1605;
  assign T1605 = T1607 ? T1606 : 12'h0;
  assign T1606 = tgts[6'hd];
  assign T1607 = hits[4'hd];
  assign T1608 = T1612 | T1609;
  assign T1609 = T1611 ? T1610 : 12'h0;
  assign T1610 = tgts[6'hc];
  assign T1611 = hits[4'hc];
  assign T1612 = T1616 | T1613;
  assign T1613 = T1615 ? T1614 : 12'h0;
  assign T1614 = tgts[6'hb];
  assign T1615 = hits[4'hb];
  assign T1616 = T1620 | T1617;
  assign T1617 = T1619 ? T1618 : 12'h0;
  assign T1618 = tgts[6'ha];
  assign T1619 = hits[4'ha];
  assign T1620 = T1624 | T1621;
  assign T1621 = T1623 ? T1622 : 12'h0;
  assign T1622 = tgts[6'h9];
  assign T1623 = hits[4'h9];
  assign T1624 = T1628 | T1625;
  assign T1625 = T1627 ? T1626 : 12'h0;
  assign T1626 = tgts[6'h8];
  assign T1627 = hits[4'h8];
  assign T1628 = T1632 | T1629;
  assign T1629 = T1631 ? T1630 : 12'h0;
  assign T1630 = tgts[6'h7];
  assign T1631 = hits[3'h7];
  assign T1632 = T1636 | T1633;
  assign T1633 = T1635 ? T1634 : 12'h0;
  assign T1634 = tgts[6'h6];
  assign T1635 = hits[3'h6];
  assign T1636 = T1640 | T1637;
  assign T1637 = T1639 ? T1638 : 12'h0;
  assign T1638 = tgts[6'h5];
  assign T1639 = hits[3'h5];
  assign T1640 = T1644 | T1641;
  assign T1641 = T1643 ? T1642 : 12'h0;
  assign T1642 = tgts[6'h4];
  assign T1643 = hits[3'h4];
  assign T1644 = T1648 | T1645;
  assign T1645 = T1647 ? T1646 : 12'h0;
  assign T1646 = tgts[6'h3];
  assign T1647 = hits[2'h3];
  assign T1648 = T1652 | T1649;
  assign T1649 = T1651 ? T1650 : 12'h0;
  assign T1650 = tgts[6'h2];
  assign T1651 = hits[2'h2];
  assign T1652 = T1656 | T1653;
  assign T1653 = T1655 ? T1654 : 12'h0;
  assign T1654 = tgts[6'h1];
  assign T1655 = hits[1'h1];
  assign T1656 = T1658 ? T1657 : 12'h0;
  assign T1657 = tgts[6'h0];
  assign T1658 = hits[1'h0];
  assign T1659 = T1848 | T1660;
  assign T1660 = T1662 ? T1661 : 27'h0;
  assign T1661 = pages[3'h5];
  assign T1662 = T1663[3'h5];
  assign T1663 = T1666 | T1664;
  assign T1664 = T1665 ? tgtPagesOH_61 : 6'h0;
  assign T1665 = hits[6'h3d];
  assign T1666 = T1669 | T1667;
  assign T1667 = T1668 ? tgtPagesOH_60 : 6'h0;
  assign T1668 = hits[6'h3c];
  assign T1669 = T1672 | T1670;
  assign T1670 = T1671 ? tgtPagesOH_59 : 6'h0;
  assign T1671 = hits[6'h3b];
  assign T1672 = T1675 | T1673;
  assign T1673 = T1674 ? tgtPagesOH_58 : 6'h0;
  assign T1674 = hits[6'h3a];
  assign T1675 = T1678 | T1676;
  assign T1676 = T1677 ? tgtPagesOH_57 : 6'h0;
  assign T1677 = hits[6'h39];
  assign T1678 = T1681 | T1679;
  assign T1679 = T1680 ? tgtPagesOH_56 : 6'h0;
  assign T1680 = hits[6'h38];
  assign T1681 = T1684 | T1682;
  assign T1682 = T1683 ? tgtPagesOH_55 : 6'h0;
  assign T1683 = hits[6'h37];
  assign T1684 = T1687 | T1685;
  assign T1685 = T1686 ? tgtPagesOH_54 : 6'h0;
  assign T1686 = hits[6'h36];
  assign T1687 = T1690 | T1688;
  assign T1688 = T1689 ? tgtPagesOH_53 : 6'h0;
  assign T1689 = hits[6'h35];
  assign T1690 = T1693 | T1691;
  assign T1691 = T1692 ? tgtPagesOH_52 : 6'h0;
  assign T1692 = hits[6'h34];
  assign T1693 = T1696 | T1694;
  assign T1694 = T1695 ? tgtPagesOH_51 : 6'h0;
  assign T1695 = hits[6'h33];
  assign T1696 = T1699 | T1697;
  assign T1697 = T1698 ? tgtPagesOH_50 : 6'h0;
  assign T1698 = hits[6'h32];
  assign T1699 = T1702 | T1700;
  assign T1700 = T1701 ? tgtPagesOH_49 : 6'h0;
  assign T1701 = hits[6'h31];
  assign T1702 = T1705 | T1703;
  assign T1703 = T1704 ? tgtPagesOH_48 : 6'h0;
  assign T1704 = hits[6'h30];
  assign T1705 = T1708 | T1706;
  assign T1706 = T1707 ? tgtPagesOH_47 : 6'h0;
  assign T1707 = hits[6'h2f];
  assign T1708 = T1711 | T1709;
  assign T1709 = T1710 ? tgtPagesOH_46 : 6'h0;
  assign T1710 = hits[6'h2e];
  assign T1711 = T1714 | T1712;
  assign T1712 = T1713 ? tgtPagesOH_45 : 6'h0;
  assign T1713 = hits[6'h2d];
  assign T1714 = T1717 | T1715;
  assign T1715 = T1716 ? tgtPagesOH_44 : 6'h0;
  assign T1716 = hits[6'h2c];
  assign T1717 = T1720 | T1718;
  assign T1718 = T1719 ? tgtPagesOH_43 : 6'h0;
  assign T1719 = hits[6'h2b];
  assign T1720 = T1723 | T1721;
  assign T1721 = T1722 ? tgtPagesOH_42 : 6'h0;
  assign T1722 = hits[6'h2a];
  assign T1723 = T1726 | T1724;
  assign T1724 = T1725 ? tgtPagesOH_41 : 6'h0;
  assign T1725 = hits[6'h29];
  assign T1726 = T1729 | T1727;
  assign T1727 = T1728 ? tgtPagesOH_40 : 6'h0;
  assign T1728 = hits[6'h28];
  assign T1729 = T1732 | T1730;
  assign T1730 = T1731 ? tgtPagesOH_39 : 6'h0;
  assign T1731 = hits[6'h27];
  assign T1732 = T1735 | T1733;
  assign T1733 = T1734 ? tgtPagesOH_38 : 6'h0;
  assign T1734 = hits[6'h26];
  assign T1735 = T1738 | T1736;
  assign T1736 = T1737 ? tgtPagesOH_37 : 6'h0;
  assign T1737 = hits[6'h25];
  assign T1738 = T1741 | T1739;
  assign T1739 = T1740 ? tgtPagesOH_36 : 6'h0;
  assign T1740 = hits[6'h24];
  assign T1741 = T1744 | T1742;
  assign T1742 = T1743 ? tgtPagesOH_35 : 6'h0;
  assign T1743 = hits[6'h23];
  assign T1744 = T1747 | T1745;
  assign T1745 = T1746 ? tgtPagesOH_34 : 6'h0;
  assign T1746 = hits[6'h22];
  assign T1747 = T1750 | T1748;
  assign T1748 = T1749 ? tgtPagesOH_33 : 6'h0;
  assign T1749 = hits[6'h21];
  assign T1750 = T1753 | T1751;
  assign T1751 = T1752 ? tgtPagesOH_32 : 6'h0;
  assign T1752 = hits[6'h20];
  assign T1753 = T1756 | T1754;
  assign T1754 = T1755 ? tgtPagesOH_31 : 6'h0;
  assign T1755 = hits[5'h1f];
  assign T1756 = T1759 | T1757;
  assign T1757 = T1758 ? tgtPagesOH_30 : 6'h0;
  assign T1758 = hits[5'h1e];
  assign T1759 = T1762 | T1760;
  assign T1760 = T1761 ? tgtPagesOH_29 : 6'h0;
  assign T1761 = hits[5'h1d];
  assign T1762 = T1765 | T1763;
  assign T1763 = T1764 ? tgtPagesOH_28 : 6'h0;
  assign T1764 = hits[5'h1c];
  assign T1765 = T1768 | T1766;
  assign T1766 = T1767 ? tgtPagesOH_27 : 6'h0;
  assign T1767 = hits[5'h1b];
  assign T1768 = T1771 | T1769;
  assign T1769 = T1770 ? tgtPagesOH_26 : 6'h0;
  assign T1770 = hits[5'h1a];
  assign T1771 = T1774 | T1772;
  assign T1772 = T1773 ? tgtPagesOH_25 : 6'h0;
  assign T1773 = hits[5'h19];
  assign T1774 = T1777 | T1775;
  assign T1775 = T1776 ? tgtPagesOH_24 : 6'h0;
  assign T1776 = hits[5'h18];
  assign T1777 = T1780 | T1778;
  assign T1778 = T1779 ? tgtPagesOH_23 : 6'h0;
  assign T1779 = hits[5'h17];
  assign T1780 = T1783 | T1781;
  assign T1781 = T1782 ? tgtPagesOH_22 : 6'h0;
  assign T1782 = hits[5'h16];
  assign T1783 = T1786 | T1784;
  assign T1784 = T1785 ? tgtPagesOH_21 : 6'h0;
  assign T1785 = hits[5'h15];
  assign T1786 = T1789 | T1787;
  assign T1787 = T1788 ? tgtPagesOH_20 : 6'h0;
  assign T1788 = hits[5'h14];
  assign T1789 = T1792 | T1790;
  assign T1790 = T1791 ? tgtPagesOH_19 : 6'h0;
  assign T1791 = hits[5'h13];
  assign T1792 = T1795 | T1793;
  assign T1793 = T1794 ? tgtPagesOH_18 : 6'h0;
  assign T1794 = hits[5'h12];
  assign T1795 = T1798 | T1796;
  assign T1796 = T1797 ? tgtPagesOH_17 : 6'h0;
  assign T1797 = hits[5'h11];
  assign T1798 = T1801 | T1799;
  assign T1799 = T1800 ? tgtPagesOH_16 : 6'h0;
  assign T1800 = hits[5'h10];
  assign T1801 = T1804 | T1802;
  assign T1802 = T1803 ? tgtPagesOH_15 : 6'h0;
  assign T1803 = hits[4'hf];
  assign T1804 = T1807 | T1805;
  assign T1805 = T1806 ? tgtPagesOH_14 : 6'h0;
  assign T1806 = hits[4'he];
  assign T1807 = T1810 | T1808;
  assign T1808 = T1809 ? tgtPagesOH_13 : 6'h0;
  assign T1809 = hits[4'hd];
  assign T1810 = T1813 | T1811;
  assign T1811 = T1812 ? tgtPagesOH_12 : 6'h0;
  assign T1812 = hits[4'hc];
  assign T1813 = T1816 | T1814;
  assign T1814 = T1815 ? tgtPagesOH_11 : 6'h0;
  assign T1815 = hits[4'hb];
  assign T1816 = T1819 | T1817;
  assign T1817 = T1818 ? tgtPagesOH_10 : 6'h0;
  assign T1818 = hits[4'ha];
  assign T1819 = T1822 | T1820;
  assign T1820 = T1821 ? tgtPagesOH_9 : 6'h0;
  assign T1821 = hits[4'h9];
  assign T1822 = T1825 | T1823;
  assign T1823 = T1824 ? tgtPagesOH_8 : 6'h0;
  assign T1824 = hits[4'h8];
  assign T1825 = T1828 | T1826;
  assign T1826 = T1827 ? tgtPagesOH_7 : 6'h0;
  assign T1827 = hits[3'h7];
  assign T1828 = T1831 | T1829;
  assign T1829 = T1830 ? tgtPagesOH_6 : 6'h0;
  assign T1830 = hits[3'h6];
  assign T1831 = T1834 | T1832;
  assign T1832 = T1833 ? tgtPagesOH_5 : 6'h0;
  assign T1833 = hits[3'h5];
  assign T1834 = T1837 | T1835;
  assign T1835 = T1836 ? tgtPagesOH_4 : 6'h0;
  assign T1836 = hits[3'h4];
  assign T1837 = T1840 | T1838;
  assign T1838 = T1839 ? tgtPagesOH_3 : 6'h0;
  assign T1839 = hits[2'h3];
  assign T1840 = T1843 | T1841;
  assign T1841 = T1842 ? tgtPagesOH_2 : 6'h0;
  assign T1842 = hits[2'h2];
  assign T1843 = T1846 | T1844;
  assign T1844 = T1845 ? tgtPagesOH_1 : 6'h0;
  assign T1845 = hits[1'h1];
  assign T1846 = T1847 ? tgtPagesOH_0 : 6'h0;
  assign T1847 = hits[1'h0];
  assign T1848 = T1852 | T1849;
  assign T1849 = T1851 ? T1850 : 27'h0;
  assign T1850 = pages[3'h4];
  assign T1851 = T1663[3'h4];
  assign T1852 = T1856 | T1853;
  assign T1853 = T1855 ? T1854 : 27'h0;
  assign T1854 = pages[3'h3];
  assign T1855 = T1663[2'h3];
  assign T1856 = T1860 | T1857;
  assign T1857 = T1859 ? T1858 : 27'h0;
  assign T1858 = pages[3'h2];
  assign T1859 = T1663[2'h2];
  assign T1860 = T1864 | T1861;
  assign T1861 = T1863 ? T1862 : 27'h0;
  assign T1862 = pages[3'h1];
  assign T1863 = T1663[1'h1];
  assign T1864 = T1866 ? T1865 : 27'h0;
  assign T1865 = pages[3'h0];
  assign T1866 = T1663[1'h0];
  assign T1867 = T1899 ? R1895 : R1868;
  assign T1869 = T1870 ? io_ras_update_bits_returnAddr : R1868;
  assign T1870 = T1894 & T1871;
  assign T1871 = T1872[1'h0];
  assign T1872 = 1'h1 << T1873;
  assign T1873 = T1874;
  assign T1874 = R1875 + 1'h1;
  assign T2348 = reset ? 1'h0 : T1876;
  assign T1876 = T1879 ? T1878 : T1877;
  assign T1877 = T1894 ? T1874 : R1875;
  assign T1878 = R1875 - 1'h1;
  assign T1879 = T1890 & T1880;
  assign T1880 = T1881 ^ 1'h1;
  assign T1881 = R1882 == 2'h0;
  assign T2349 = reset ? 2'h0 : T1883;
  assign T1883 = io_invalidate ? 2'h0 : T1884;
  assign T1884 = T1879 ? T1889 : T1885;
  assign T1885 = T1887 ? T1886 : R1882;
  assign T1886 = R1882 + 2'h1;
  assign T1887 = T1894 & T1888;
  assign T1888 = R1882 < 2'h2;
  assign T1889 = R1882 - 2'h1;
  assign T1890 = io_ras_update_valid & T1891;
  assign T1891 = T1893 & T1892;
  assign T1892 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T1893 = io_ras_update_bits_isCall ^ 1'h1;
  assign T1894 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T1896 = T1897 ? io_ras_update_bits_returnAddr : R1895;
  assign T1897 = T1894 & T1898;
  assign T1898 = T1872[1'h1];
  assign T1899 = R1875;
  assign T1900 = T2276 & T1901;
  assign T1901 = T1911 | T1902;
  assign T1902 = T1910 ? useRAS_61 : 1'h0;
  assign T1903 = T1906 ? R1904 : useRAS_61;
  assign T1905 = io_btb_update_valid ? io_btb_update_bits_isReturn : R1904;
  assign T1906 = R7 & T1907;
  assign T1907 = T1908[6'h3d];
  assign T1908 = 1'h1 << T1909;
  assign T1909 = T42;
  assign T1910 = hits[6'h3d];
  assign T1911 = T1917 | T1912;
  assign T1912 = T1916 ? useRAS_60 : 1'h0;
  assign T1913 = T1914 ? R1904 : useRAS_60;
  assign T1914 = R7 & T1915;
  assign T1915 = T1908[6'h3c];
  assign T1916 = hits[6'h3c];
  assign T1917 = T1923 | T1918;
  assign T1918 = T1922 ? useRAS_59 : 1'h0;
  assign T1919 = T1920 ? R1904 : useRAS_59;
  assign T1920 = R7 & T1921;
  assign T1921 = T1908[6'h3b];
  assign T1922 = hits[6'h3b];
  assign T1923 = T1929 | T1924;
  assign T1924 = T1928 ? useRAS_58 : 1'h0;
  assign T1925 = T1926 ? R1904 : useRAS_58;
  assign T1926 = R7 & T1927;
  assign T1927 = T1908[6'h3a];
  assign T1928 = hits[6'h3a];
  assign T1929 = T1935 | T1930;
  assign T1930 = T1934 ? useRAS_57 : 1'h0;
  assign T1931 = T1932 ? R1904 : useRAS_57;
  assign T1932 = R7 & T1933;
  assign T1933 = T1908[6'h39];
  assign T1934 = hits[6'h39];
  assign T1935 = T1941 | T1936;
  assign T1936 = T1940 ? useRAS_56 : 1'h0;
  assign T1937 = T1938 ? R1904 : useRAS_56;
  assign T1938 = R7 & T1939;
  assign T1939 = T1908[6'h38];
  assign T1940 = hits[6'h38];
  assign T1941 = T1947 | T1942;
  assign T1942 = T1946 ? useRAS_55 : 1'h0;
  assign T1943 = T1944 ? R1904 : useRAS_55;
  assign T1944 = R7 & T1945;
  assign T1945 = T1908[6'h37];
  assign T1946 = hits[6'h37];
  assign T1947 = T1953 | T1948;
  assign T1948 = T1952 ? useRAS_54 : 1'h0;
  assign T1949 = T1950 ? R1904 : useRAS_54;
  assign T1950 = R7 & T1951;
  assign T1951 = T1908[6'h36];
  assign T1952 = hits[6'h36];
  assign T1953 = T1959 | T1954;
  assign T1954 = T1958 ? useRAS_53 : 1'h0;
  assign T1955 = T1956 ? R1904 : useRAS_53;
  assign T1956 = R7 & T1957;
  assign T1957 = T1908[6'h35];
  assign T1958 = hits[6'h35];
  assign T1959 = T1965 | T1960;
  assign T1960 = T1964 ? useRAS_52 : 1'h0;
  assign T1961 = T1962 ? R1904 : useRAS_52;
  assign T1962 = R7 & T1963;
  assign T1963 = T1908[6'h34];
  assign T1964 = hits[6'h34];
  assign T1965 = T1971 | T1966;
  assign T1966 = T1970 ? useRAS_51 : 1'h0;
  assign T1967 = T1968 ? R1904 : useRAS_51;
  assign T1968 = R7 & T1969;
  assign T1969 = T1908[6'h33];
  assign T1970 = hits[6'h33];
  assign T1971 = T1977 | T1972;
  assign T1972 = T1976 ? useRAS_50 : 1'h0;
  assign T1973 = T1974 ? R1904 : useRAS_50;
  assign T1974 = R7 & T1975;
  assign T1975 = T1908[6'h32];
  assign T1976 = hits[6'h32];
  assign T1977 = T1983 | T1978;
  assign T1978 = T1982 ? useRAS_49 : 1'h0;
  assign T1979 = T1980 ? R1904 : useRAS_49;
  assign T1980 = R7 & T1981;
  assign T1981 = T1908[6'h31];
  assign T1982 = hits[6'h31];
  assign T1983 = T1989 | T1984;
  assign T1984 = T1988 ? useRAS_48 : 1'h0;
  assign T1985 = T1986 ? R1904 : useRAS_48;
  assign T1986 = R7 & T1987;
  assign T1987 = T1908[6'h30];
  assign T1988 = hits[6'h30];
  assign T1989 = T1995 | T1990;
  assign T1990 = T1994 ? useRAS_47 : 1'h0;
  assign T1991 = T1992 ? R1904 : useRAS_47;
  assign T1992 = R7 & T1993;
  assign T1993 = T1908[6'h2f];
  assign T1994 = hits[6'h2f];
  assign T1995 = T2001 | T1996;
  assign T1996 = T2000 ? useRAS_46 : 1'h0;
  assign T1997 = T1998 ? R1904 : useRAS_46;
  assign T1998 = R7 & T1999;
  assign T1999 = T1908[6'h2e];
  assign T2000 = hits[6'h2e];
  assign T2001 = T2007 | T2002;
  assign T2002 = T2006 ? useRAS_45 : 1'h0;
  assign T2003 = T2004 ? R1904 : useRAS_45;
  assign T2004 = R7 & T2005;
  assign T2005 = T1908[6'h2d];
  assign T2006 = hits[6'h2d];
  assign T2007 = T2013 | T2008;
  assign T2008 = T2012 ? useRAS_44 : 1'h0;
  assign T2009 = T2010 ? R1904 : useRAS_44;
  assign T2010 = R7 & T2011;
  assign T2011 = T1908[6'h2c];
  assign T2012 = hits[6'h2c];
  assign T2013 = T2019 | T2014;
  assign T2014 = T2018 ? useRAS_43 : 1'h0;
  assign T2015 = T2016 ? R1904 : useRAS_43;
  assign T2016 = R7 & T2017;
  assign T2017 = T1908[6'h2b];
  assign T2018 = hits[6'h2b];
  assign T2019 = T2025 | T2020;
  assign T2020 = T2024 ? useRAS_42 : 1'h0;
  assign T2021 = T2022 ? R1904 : useRAS_42;
  assign T2022 = R7 & T2023;
  assign T2023 = T1908[6'h2a];
  assign T2024 = hits[6'h2a];
  assign T2025 = T2031 | T2026;
  assign T2026 = T2030 ? useRAS_41 : 1'h0;
  assign T2027 = T2028 ? R1904 : useRAS_41;
  assign T2028 = R7 & T2029;
  assign T2029 = T1908[6'h29];
  assign T2030 = hits[6'h29];
  assign T2031 = T2037 | T2032;
  assign T2032 = T2036 ? useRAS_40 : 1'h0;
  assign T2033 = T2034 ? R1904 : useRAS_40;
  assign T2034 = R7 & T2035;
  assign T2035 = T1908[6'h28];
  assign T2036 = hits[6'h28];
  assign T2037 = T2043 | T2038;
  assign T2038 = T2042 ? useRAS_39 : 1'h0;
  assign T2039 = T2040 ? R1904 : useRAS_39;
  assign T2040 = R7 & T2041;
  assign T2041 = T1908[6'h27];
  assign T2042 = hits[6'h27];
  assign T2043 = T2049 | T2044;
  assign T2044 = T2048 ? useRAS_38 : 1'h0;
  assign T2045 = T2046 ? R1904 : useRAS_38;
  assign T2046 = R7 & T2047;
  assign T2047 = T1908[6'h26];
  assign T2048 = hits[6'h26];
  assign T2049 = T2055 | T2050;
  assign T2050 = T2054 ? useRAS_37 : 1'h0;
  assign T2051 = T2052 ? R1904 : useRAS_37;
  assign T2052 = R7 & T2053;
  assign T2053 = T1908[6'h25];
  assign T2054 = hits[6'h25];
  assign T2055 = T2061 | T2056;
  assign T2056 = T2060 ? useRAS_36 : 1'h0;
  assign T2057 = T2058 ? R1904 : useRAS_36;
  assign T2058 = R7 & T2059;
  assign T2059 = T1908[6'h24];
  assign T2060 = hits[6'h24];
  assign T2061 = T2067 | T2062;
  assign T2062 = T2066 ? useRAS_35 : 1'h0;
  assign T2063 = T2064 ? R1904 : useRAS_35;
  assign T2064 = R7 & T2065;
  assign T2065 = T1908[6'h23];
  assign T2066 = hits[6'h23];
  assign T2067 = T2073 | T2068;
  assign T2068 = T2072 ? useRAS_34 : 1'h0;
  assign T2069 = T2070 ? R1904 : useRAS_34;
  assign T2070 = R7 & T2071;
  assign T2071 = T1908[6'h22];
  assign T2072 = hits[6'h22];
  assign T2073 = T2079 | T2074;
  assign T2074 = T2078 ? useRAS_33 : 1'h0;
  assign T2075 = T2076 ? R1904 : useRAS_33;
  assign T2076 = R7 & T2077;
  assign T2077 = T1908[6'h21];
  assign T2078 = hits[6'h21];
  assign T2079 = T2085 | T2080;
  assign T2080 = T2084 ? useRAS_32 : 1'h0;
  assign T2081 = T2082 ? R1904 : useRAS_32;
  assign T2082 = R7 & T2083;
  assign T2083 = T1908[6'h20];
  assign T2084 = hits[6'h20];
  assign T2085 = T2091 | T2086;
  assign T2086 = T2090 ? useRAS_31 : 1'h0;
  assign T2087 = T2088 ? R1904 : useRAS_31;
  assign T2088 = R7 & T2089;
  assign T2089 = T1908[5'h1f];
  assign T2090 = hits[5'h1f];
  assign T2091 = T2097 | T2092;
  assign T2092 = T2096 ? useRAS_30 : 1'h0;
  assign T2093 = T2094 ? R1904 : useRAS_30;
  assign T2094 = R7 & T2095;
  assign T2095 = T1908[5'h1e];
  assign T2096 = hits[5'h1e];
  assign T2097 = T2103 | T2098;
  assign T2098 = T2102 ? useRAS_29 : 1'h0;
  assign T2099 = T2100 ? R1904 : useRAS_29;
  assign T2100 = R7 & T2101;
  assign T2101 = T1908[5'h1d];
  assign T2102 = hits[5'h1d];
  assign T2103 = T2109 | T2104;
  assign T2104 = T2108 ? useRAS_28 : 1'h0;
  assign T2105 = T2106 ? R1904 : useRAS_28;
  assign T2106 = R7 & T2107;
  assign T2107 = T1908[5'h1c];
  assign T2108 = hits[5'h1c];
  assign T2109 = T2115 | T2110;
  assign T2110 = T2114 ? useRAS_27 : 1'h0;
  assign T2111 = T2112 ? R1904 : useRAS_27;
  assign T2112 = R7 & T2113;
  assign T2113 = T1908[5'h1b];
  assign T2114 = hits[5'h1b];
  assign T2115 = T2121 | T2116;
  assign T2116 = T2120 ? useRAS_26 : 1'h0;
  assign T2117 = T2118 ? R1904 : useRAS_26;
  assign T2118 = R7 & T2119;
  assign T2119 = T1908[5'h1a];
  assign T2120 = hits[5'h1a];
  assign T2121 = T2127 | T2122;
  assign T2122 = T2126 ? useRAS_25 : 1'h0;
  assign T2123 = T2124 ? R1904 : useRAS_25;
  assign T2124 = R7 & T2125;
  assign T2125 = T1908[5'h19];
  assign T2126 = hits[5'h19];
  assign T2127 = T2133 | T2128;
  assign T2128 = T2132 ? useRAS_24 : 1'h0;
  assign T2129 = T2130 ? R1904 : useRAS_24;
  assign T2130 = R7 & T2131;
  assign T2131 = T1908[5'h18];
  assign T2132 = hits[5'h18];
  assign T2133 = T2139 | T2134;
  assign T2134 = T2138 ? useRAS_23 : 1'h0;
  assign T2135 = T2136 ? R1904 : useRAS_23;
  assign T2136 = R7 & T2137;
  assign T2137 = T1908[5'h17];
  assign T2138 = hits[5'h17];
  assign T2139 = T2145 | T2140;
  assign T2140 = T2144 ? useRAS_22 : 1'h0;
  assign T2141 = T2142 ? R1904 : useRAS_22;
  assign T2142 = R7 & T2143;
  assign T2143 = T1908[5'h16];
  assign T2144 = hits[5'h16];
  assign T2145 = T2151 | T2146;
  assign T2146 = T2150 ? useRAS_21 : 1'h0;
  assign T2147 = T2148 ? R1904 : useRAS_21;
  assign T2148 = R7 & T2149;
  assign T2149 = T1908[5'h15];
  assign T2150 = hits[5'h15];
  assign T2151 = T2157 | T2152;
  assign T2152 = T2156 ? useRAS_20 : 1'h0;
  assign T2153 = T2154 ? R1904 : useRAS_20;
  assign T2154 = R7 & T2155;
  assign T2155 = T1908[5'h14];
  assign T2156 = hits[5'h14];
  assign T2157 = T2163 | T2158;
  assign T2158 = T2162 ? useRAS_19 : 1'h0;
  assign T2159 = T2160 ? R1904 : useRAS_19;
  assign T2160 = R7 & T2161;
  assign T2161 = T1908[5'h13];
  assign T2162 = hits[5'h13];
  assign T2163 = T2169 | T2164;
  assign T2164 = T2168 ? useRAS_18 : 1'h0;
  assign T2165 = T2166 ? R1904 : useRAS_18;
  assign T2166 = R7 & T2167;
  assign T2167 = T1908[5'h12];
  assign T2168 = hits[5'h12];
  assign T2169 = T2175 | T2170;
  assign T2170 = T2174 ? useRAS_17 : 1'h0;
  assign T2171 = T2172 ? R1904 : useRAS_17;
  assign T2172 = R7 & T2173;
  assign T2173 = T1908[5'h11];
  assign T2174 = hits[5'h11];
  assign T2175 = T2181 | T2176;
  assign T2176 = T2180 ? useRAS_16 : 1'h0;
  assign T2177 = T2178 ? R1904 : useRAS_16;
  assign T2178 = R7 & T2179;
  assign T2179 = T1908[5'h10];
  assign T2180 = hits[5'h10];
  assign T2181 = T2187 | T2182;
  assign T2182 = T2186 ? useRAS_15 : 1'h0;
  assign T2183 = T2184 ? R1904 : useRAS_15;
  assign T2184 = R7 & T2185;
  assign T2185 = T1908[4'hf];
  assign T2186 = hits[4'hf];
  assign T2187 = T2193 | T2188;
  assign T2188 = T2192 ? useRAS_14 : 1'h0;
  assign T2189 = T2190 ? R1904 : useRAS_14;
  assign T2190 = R7 & T2191;
  assign T2191 = T1908[4'he];
  assign T2192 = hits[4'he];
  assign T2193 = T2199 | T2194;
  assign T2194 = T2198 ? useRAS_13 : 1'h0;
  assign T2195 = T2196 ? R1904 : useRAS_13;
  assign T2196 = R7 & T2197;
  assign T2197 = T1908[4'hd];
  assign T2198 = hits[4'hd];
  assign T2199 = T2205 | T2200;
  assign T2200 = T2204 ? useRAS_12 : 1'h0;
  assign T2201 = T2202 ? R1904 : useRAS_12;
  assign T2202 = R7 & T2203;
  assign T2203 = T1908[4'hc];
  assign T2204 = hits[4'hc];
  assign T2205 = T2211 | T2206;
  assign T2206 = T2210 ? useRAS_11 : 1'h0;
  assign T2207 = T2208 ? R1904 : useRAS_11;
  assign T2208 = R7 & T2209;
  assign T2209 = T1908[4'hb];
  assign T2210 = hits[4'hb];
  assign T2211 = T2217 | T2212;
  assign T2212 = T2216 ? useRAS_10 : 1'h0;
  assign T2213 = T2214 ? R1904 : useRAS_10;
  assign T2214 = R7 & T2215;
  assign T2215 = T1908[4'ha];
  assign T2216 = hits[4'ha];
  assign T2217 = T2223 | T2218;
  assign T2218 = T2222 ? useRAS_9 : 1'h0;
  assign T2219 = T2220 ? R1904 : useRAS_9;
  assign T2220 = R7 & T2221;
  assign T2221 = T1908[4'h9];
  assign T2222 = hits[4'h9];
  assign T2223 = T2229 | T2224;
  assign T2224 = T2228 ? useRAS_8 : 1'h0;
  assign T2225 = T2226 ? R1904 : useRAS_8;
  assign T2226 = R7 & T2227;
  assign T2227 = T1908[4'h8];
  assign T2228 = hits[4'h8];
  assign T2229 = T2235 | T2230;
  assign T2230 = T2234 ? useRAS_7 : 1'h0;
  assign T2231 = T2232 ? R1904 : useRAS_7;
  assign T2232 = R7 & T2233;
  assign T2233 = T1908[3'h7];
  assign T2234 = hits[3'h7];
  assign T2235 = T2241 | T2236;
  assign T2236 = T2240 ? useRAS_6 : 1'h0;
  assign T2237 = T2238 ? R1904 : useRAS_6;
  assign T2238 = R7 & T2239;
  assign T2239 = T1908[3'h6];
  assign T2240 = hits[3'h6];
  assign T2241 = T2247 | T2242;
  assign T2242 = T2246 ? useRAS_5 : 1'h0;
  assign T2243 = T2244 ? R1904 : useRAS_5;
  assign T2244 = R7 & T2245;
  assign T2245 = T1908[3'h5];
  assign T2246 = hits[3'h5];
  assign T2247 = T2253 | T2248;
  assign T2248 = T2252 ? useRAS_4 : 1'h0;
  assign T2249 = T2250 ? R1904 : useRAS_4;
  assign T2250 = R7 & T2251;
  assign T2251 = T1908[3'h4];
  assign T2252 = hits[3'h4];
  assign T2253 = T2259 | T2254;
  assign T2254 = T2258 ? useRAS_3 : 1'h0;
  assign T2255 = T2256 ? R1904 : useRAS_3;
  assign T2256 = R7 & T2257;
  assign T2257 = T1908[2'h3];
  assign T2258 = hits[2'h3];
  assign T2259 = T2265 | T2260;
  assign T2260 = T2264 ? useRAS_2 : 1'h0;
  assign T2261 = T2262 ? R1904 : useRAS_2;
  assign T2262 = R7 & T2263;
  assign T2263 = T1908[2'h2];
  assign T2264 = hits[2'h2];
  assign T2265 = T2271 | T2266;
  assign T2266 = T2270 ? useRAS_1 : 1'h0;
  assign T2267 = T2268 ? R1904 : useRAS_1;
  assign T2268 = R7 & T2269;
  assign T2269 = T1908[1'h1];
  assign T2270 = hits[1'h1];
  assign T2271 = T2275 ? useRAS_0 : 1'h0;
  assign T2272 = T2273 ? R1904 : useRAS_0;
  assign T2273 = R7 & T2274;
  assign T2274 = T1908[1'h0];
  assign T2275 = hits[1'h0];
  assign T2276 = T2277 ^ 1'h1;
  assign T2277 = R1882 == 2'h0;
  assign T2278 = T1894 & T1901;
  assign io_resp_bits_bridx = T2279;
  assign T2279 = brIdx[io_resp_bits_entry];
  assign T2281 = R7 & T2282;
  assign T2282 = T42 < 6'h3e;
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_taken = T2283;
  assign T2283 = T2284 ? 1'h0 : io_resp_valid;
  assign T2284 = T2285 & T32;
  assign T2285 = T2286 ^ 1'h1;
  assign T2286 = T8[1'h0];
  assign io_resp_valid = T2287;
  assign T2287 = hits != 62'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
// synthesis translate_on
`endif
    if(io_btb_update_valid) begin
      R4 <= io_btb_update_bits_target;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_btb_update_valid;
    end
    if (T21)
      T10[T22] <= T12;
    if(T1402) begin
      R25 <= T1400;
    end else if(T31) begin
      R25 <= T28;
    end
    if(T38) begin
      isJump_61 <= R36;
    end
    if(io_btb_update_valid) begin
      R36 <= io_btb_update_bits_isJump;
    end
    if(reset) begin
      nextRepl <= 6'h0;
    end else if(T47) begin
      nextRepl <= T44;
    end
    if(io_btb_update_valid) begin
      R49 <= io_btb_update_bits_prediction_bits_entry;
    end
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end
    if(reset) begin
      pageValid <= 6'h0;
    end else if(io_invalidate) begin
      pageValid <= 6'h0;
    end else if(T137) begin
      pageValid <= T64;
    end
    if(reset) begin
      R70 <= 3'h0;
    end else if(T75) begin
      R70 <= T72;
    end
    if(io_btb_update_valid) begin
      R82 <= io_btb_update_bits_pc;
    end
    if (T91)
      pages[3'h5] <= T86;
    if (T96)
      pages[3'h3] <= T86;
    if (T100)
      pages[3'h1] <= T86;
    if (T107)
      pages[3'h4] <= T104;
    if (T112)
      pages[3'h2] <= T104;
    if (T116)
      pages[3'h0] <= T104;
    if (T160)
      idxPages[T42] <= T2294;
    if (T473)
      idxs[T42] <= T2305;
    idxValid <= T2306;
    if (T672)
      tgtPages[T42] <= T2310;
    if(T1037) begin
      isJump_60 <= R36;
    end
    if(T1043) begin
      isJump_59 <= R36;
    end
    if(T1049) begin
      isJump_58 <= R36;
    end
    if(T1055) begin
      isJump_57 <= R36;
    end
    if(T1061) begin
      isJump_56 <= R36;
    end
    if(T1067) begin
      isJump_55 <= R36;
    end
    if(T1073) begin
      isJump_54 <= R36;
    end
    if(T1079) begin
      isJump_53 <= R36;
    end
    if(T1085) begin
      isJump_52 <= R36;
    end
    if(T1091) begin
      isJump_51 <= R36;
    end
    if(T1097) begin
      isJump_50 <= R36;
    end
    if(T1103) begin
      isJump_49 <= R36;
    end
    if(T1109) begin
      isJump_48 <= R36;
    end
    if(T1115) begin
      isJump_47 <= R36;
    end
    if(T1121) begin
      isJump_46 <= R36;
    end
    if(T1127) begin
      isJump_45 <= R36;
    end
    if(T1133) begin
      isJump_44 <= R36;
    end
    if(T1139) begin
      isJump_43 <= R36;
    end
    if(T1145) begin
      isJump_42 <= R36;
    end
    if(T1151) begin
      isJump_41 <= R36;
    end
    if(T1157) begin
      isJump_40 <= R36;
    end
    if(T1163) begin
      isJump_39 <= R36;
    end
    if(T1169) begin
      isJump_38 <= R36;
    end
    if(T1175) begin
      isJump_37 <= R36;
    end
    if(T1181) begin
      isJump_36 <= R36;
    end
    if(T1187) begin
      isJump_35 <= R36;
    end
    if(T1193) begin
      isJump_34 <= R36;
    end
    if(T1199) begin
      isJump_33 <= R36;
    end
    if(T1205) begin
      isJump_32 <= R36;
    end
    if(T1211) begin
      isJump_31 <= R36;
    end
    if(T1217) begin
      isJump_30 <= R36;
    end
    if(T1223) begin
      isJump_29 <= R36;
    end
    if(T1229) begin
      isJump_28 <= R36;
    end
    if(T1235) begin
      isJump_27 <= R36;
    end
    if(T1241) begin
      isJump_26 <= R36;
    end
    if(T1247) begin
      isJump_25 <= R36;
    end
    if(T1253) begin
      isJump_24 <= R36;
    end
    if(T1259) begin
      isJump_23 <= R36;
    end
    if(T1265) begin
      isJump_22 <= R36;
    end
    if(T1271) begin
      isJump_21 <= R36;
    end
    if(T1277) begin
      isJump_20 <= R36;
    end
    if(T1283) begin
      isJump_19 <= R36;
    end
    if(T1289) begin
      isJump_18 <= R36;
    end
    if(T1295) begin
      isJump_17 <= R36;
    end
    if(T1301) begin
      isJump_16 <= R36;
    end
    if(T1307) begin
      isJump_15 <= R36;
    end
    if(T1313) begin
      isJump_14 <= R36;
    end
    if(T1319) begin
      isJump_13 <= R36;
    end
    if(T1325) begin
      isJump_12 <= R36;
    end
    if(T1331) begin
      isJump_11 <= R36;
    end
    if(T1337) begin
      isJump_10 <= R36;
    end
    if(T1343) begin
      isJump_9 <= R36;
    end
    if(T1349) begin
      isJump_8 <= R36;
    end
    if(T1355) begin
      isJump_7 <= R36;
    end
    if(T1361) begin
      isJump_6 <= R36;
    end
    if(T1367) begin
      isJump_5 <= R36;
    end
    if(T1373) begin
      isJump_4 <= R36;
    end
    if(T1379) begin
      isJump_3 <= R36;
    end
    if(T1385) begin
      isJump_2 <= R36;
    end
    if(T1391) begin
      isJump_1 <= R36;
    end
    if(T1396) begin
      isJump_0 <= R36;
    end
    if (T1413)
      tgts[T42] <= T2347;
    if(T1870) begin
      R1868 <= io_ras_update_bits_returnAddr;
    end
    if(reset) begin
      R1875 <= 1'h0;
    end else if(T1879) begin
      R1875 <= T1878;
    end else if(T1894) begin
      R1875 <= T1874;
    end
    if(reset) begin
      R1882 <= 2'h0;
    end else if(io_invalidate) begin
      R1882 <= 2'h0;
    end else if(T1879) begin
      R1882 <= T1889;
    end else if(T1887) begin
      R1882 <= T1886;
    end
    if(T1897) begin
      R1895 <= io_ras_update_bits_returnAddr;
    end
    if(T1906) begin
      useRAS_61 <= R1904;
    end
    if(io_btb_update_valid) begin
      R1904 <= io_btb_update_bits_isReturn;
    end
    if(T1914) begin
      useRAS_60 <= R1904;
    end
    if(T1920) begin
      useRAS_59 <= R1904;
    end
    if(T1926) begin
      useRAS_58 <= R1904;
    end
    if(T1932) begin
      useRAS_57 <= R1904;
    end
    if(T1938) begin
      useRAS_56 <= R1904;
    end
    if(T1944) begin
      useRAS_55 <= R1904;
    end
    if(T1950) begin
      useRAS_54 <= R1904;
    end
    if(T1956) begin
      useRAS_53 <= R1904;
    end
    if(T1962) begin
      useRAS_52 <= R1904;
    end
    if(T1968) begin
      useRAS_51 <= R1904;
    end
    if(T1974) begin
      useRAS_50 <= R1904;
    end
    if(T1980) begin
      useRAS_49 <= R1904;
    end
    if(T1986) begin
      useRAS_48 <= R1904;
    end
    if(T1992) begin
      useRAS_47 <= R1904;
    end
    if(T1998) begin
      useRAS_46 <= R1904;
    end
    if(T2004) begin
      useRAS_45 <= R1904;
    end
    if(T2010) begin
      useRAS_44 <= R1904;
    end
    if(T2016) begin
      useRAS_43 <= R1904;
    end
    if(T2022) begin
      useRAS_42 <= R1904;
    end
    if(T2028) begin
      useRAS_41 <= R1904;
    end
    if(T2034) begin
      useRAS_40 <= R1904;
    end
    if(T2040) begin
      useRAS_39 <= R1904;
    end
    if(T2046) begin
      useRAS_38 <= R1904;
    end
    if(T2052) begin
      useRAS_37 <= R1904;
    end
    if(T2058) begin
      useRAS_36 <= R1904;
    end
    if(T2064) begin
      useRAS_35 <= R1904;
    end
    if(T2070) begin
      useRAS_34 <= R1904;
    end
    if(T2076) begin
      useRAS_33 <= R1904;
    end
    if(T2082) begin
      useRAS_32 <= R1904;
    end
    if(T2088) begin
      useRAS_31 <= R1904;
    end
    if(T2094) begin
      useRAS_30 <= R1904;
    end
    if(T2100) begin
      useRAS_29 <= R1904;
    end
    if(T2106) begin
      useRAS_28 <= R1904;
    end
    if(T2112) begin
      useRAS_27 <= R1904;
    end
    if(T2118) begin
      useRAS_26 <= R1904;
    end
    if(T2124) begin
      useRAS_25 <= R1904;
    end
    if(T2130) begin
      useRAS_24 <= R1904;
    end
    if(T2136) begin
      useRAS_23 <= R1904;
    end
    if(T2142) begin
      useRAS_22 <= R1904;
    end
    if(T2148) begin
      useRAS_21 <= R1904;
    end
    if(T2154) begin
      useRAS_20 <= R1904;
    end
    if(T2160) begin
      useRAS_19 <= R1904;
    end
    if(T2166) begin
      useRAS_18 <= R1904;
    end
    if(T2172) begin
      useRAS_17 <= R1904;
    end
    if(T2178) begin
      useRAS_16 <= R1904;
    end
    if(T2184) begin
      useRAS_15 <= R1904;
    end
    if(T2190) begin
      useRAS_14 <= R1904;
    end
    if(T2196) begin
      useRAS_13 <= R1904;
    end
    if(T2202) begin
      useRAS_12 <= R1904;
    end
    if(T2208) begin
      useRAS_11 <= R1904;
    end
    if(T2214) begin
      useRAS_10 <= R1904;
    end
    if(T2220) begin
      useRAS_9 <= R1904;
    end
    if(T2226) begin
      useRAS_8 <= R1904;
    end
    if(T2232) begin
      useRAS_7 <= R1904;
    end
    if(T2238) begin
      useRAS_6 <= R1904;
    end
    if(T2244) begin
      useRAS_5 <= R1904;
    end
    if(T2250) begin
      useRAS_4 <= R1904;
    end
    if(T2256) begin
      useRAS_3 <= R1904;
    end
    if(T2262) begin
      useRAS_2 <= R1904;
    end
    if(T2268) begin
      useRAS_1 <= R1904;
    end
    if(T2273) begin
      useRAS_0 <= R1904;
    end
    if (T2281)
      brIdx[T42] <= 1'h0;
  end
endmodule

module FlowThroughSerializer(
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_addr_beat,
    input [5:0] io_in_bits_client_xact_id,
    input [3:0] io_in_bits_manager_xact_id,
    input  io_in_bits_is_builtin_type,
    input [3:0] io_in_bits_g_type,
    input [127:0] io_in_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[5:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output io_cnt,
    output io_done
);



  assign io_done = 1'h1;
  assign io_cnt = 1'h0;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_valid = io_in_valid;
  assign io_in_ready = io_out_ready;
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [11:0] io_req_bits_idx,
    input [19:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    //output[31:0] io_resp_bits_data
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[5:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  init
);

  wire[127:0] T0;
  wire[16:0] T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[5:0] T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] refill_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [11:0] s1_pgoff;
  wire[11:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s1_miss;
  wire T14;
  wire s1_any_tag_hit;
  wire T15;
  wire T16;
  wire T17;
  wire s1_disparity_3;
  wire T18;
  wire s1_disparity_2;
  wire T19;
  wire s1_disparity_1;
  wire s1_disparity_0;
  wire T20;
  wire s1_tag_hit_3;
  wire T21;
  wire s1_tag_match_3;
  wire T22;
  wire[19:0] s1_tag;
  wire[19:0] T23;
  wire[79:0] T24;
  wire T80;
  wire s0_valid;
  wire T81;
  wire stall;
  reg  s1_valid;
  wire T230;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T82;
  wire refill_done;
  wire refill_wrap;
  wire T54;
  reg [1:0] refill_cnt;
  wire[1:0] T231;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  reg [1:0] state;
  wire[1:0] T232;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[5:0] T73;
  wire[11:0] s0_pgoff;
  wire T74;
  wire[79:0] T25;
  wire[79:0] T26;
  wire[79:0] T27;
  wire[39:0] T28;
  wire[19:0] T29;
  wire[19:0] T233;
  wire T30;
  wire[1:0] repl_way;
  reg [15:0] R31;
  wire[15:0] T234;
  wire[15:0] T32;
  wire[15:0] T33;
  wire[14:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[19:0] T42;
  wire[19:0] T235;
  wire T43;
  wire[39:0] T44;
  wire[19:0] T45;
  wire[19:0] T236;
  wire T46;
  wire[19:0] T47;
  wire[19:0] T237;
  wire T48;
  wire[79:0] T49;
  wire[79:0] T50;
  wire[39:0] T51;
  wire[19:0] T52;
  wire[19:0] refill_tag;
  wire[39:0] T53;
  wire[5:0] s1_idx;
  reg [5:0] R71;
  wire[5:0] T72;
  wire T83;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire[5:0] T87;
  reg [255:0] vb_array;
  wire[255:0] T238;
  wire[255:0] T88;
  wire[255:0] T89;
  wire[255:0] T90;
  wire[255:0] T91;
  wire[255:0] T92;
  wire[255:0] T93;
  wire[255:0] T94;
  wire[255:0] T95;
  wire[255:0] T96;
  wire[7:0] T97;
  wire[255:0] T239;
  wire T98;
  wire[255:0] T99;
  wire[255:0] T100;
  wire T101;
  wire T102;
  reg  invalidated;
  wire T103;
  wire T104;
  wire[255:0] T105;
  wire[255:0] T240;
  wire[127:0] T106;
  wire[127:0] T107;
  wire[6:0] T108;
  wire[127:0] T241;
  wire T109;
  wire[127:0] T242;
  wire T243;
  wire[255:0] T110;
  wire[255:0] T244;
  wire[127:0] T111;
  wire T112;
  wire[255:0] T113;
  wire[255:0] T245;
  wire[127:0] T114;
  wire[127:0] T115;
  wire[6:0] T116;
  wire[127:0] T246;
  wire T117;
  wire[127:0] T247;
  wire T248;
  wire[255:0] T118;
  wire[255:0] T249;
  wire[127:0] T119;
  wire T120;
  wire[255:0] T121;
  wire[255:0] T122;
  wire[255:0] T123;
  wire[7:0] T124;
  wire[255:0] T250;
  wire T125;
  wire[255:0] T126;
  wire[255:0] T127;
  wire T128;
  wire[255:0] T129;
  wire[255:0] T130;
  wire[255:0] T131;
  wire[7:0] T132;
  wire[255:0] T251;
  wire T133;
  wire[255:0] T134;
  wire[255:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire s1_tag_hit_2;
  wire T139;
  wire s1_tag_match_2;
  wire T140;
  wire[19:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[7:0] T145;
  wire[5:0] T146;
  wire T147;
  wire T148;
  wire s1_tag_hit_1;
  wire T149;
  wire s1_tag_match_1;
  wire T150;
  wire[19:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire[6:0] T155;
  wire[5:0] T156;
  wire T157;
  wire s1_tag_hit_0;
  wire T158;
  wire s1_tag_match_0;
  wire T159;
  wire[19:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire[6:0] T164;
  wire[5:0] T165;
  wire T166;
  wire out_valid;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[127:0] T175;
  wire[127:0] T176;
  wire[127:0] s1_dout_3;
  wire[127:0] T177;
  wire T187;
  wire T188;
  wire T181;
  wire T182;
  wire[7:0] T186;
  wire[127:0] T179;
  wire[127:0] T180;
  wire[7:0] T183;
  reg [7:0] R184;
  wire[7:0] T185;
  wire[127:0] T189;
  wire[127:0] T190;
  wire[127:0] s1_dout_2;
  wire[127:0] T191;
  wire T201;
  wire T202;
  wire T195;
  wire T196;
  wire[7:0] T200;
  wire[127:0] T193;
  wire[127:0] T194;
  wire[7:0] T197;
  reg [7:0] R198;
  wire[7:0] T199;
  wire[127:0] T203;
  wire[127:0] T204;
  wire[127:0] s1_dout_1;
  wire[127:0] T205;
  wire T215;
  wire T216;
  wire T209;
  wire T210;
  wire[7:0] T214;
  wire[127:0] T207;
  wire[127:0] T208;
  wire[7:0] T211;
  reg [7:0] R212;
  wire[7:0] T213;
  wire[127:0] T217;
  wire[127:0] s1_dout_0;
  wire[127:0] T218;
  wire T228;
  wire T229;
  wire T222;
  wire T223;
  wire[7:0] T227;
  wire[127:0] T220;
  wire[127:0] T221;
  wire[7:0] T224;
  reg [7:0] R225;
  wire[7:0] T226;
  wire s1_hit;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    refill_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    s1_valid = {1{$random}};
    refill_cnt = {1{$random}};
    state = {1{$random}};
    R31 = {1{$random}};
    R71 = {1{$random}};
    vb_array = {8{$random}};
    invalidated = {1{$random}};
    R184 = {1{$random}};
    R198 = {1{$random}};
    R212 = {1{$random}};
    R225 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_resp_bits_data = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = T0;
  assign T0 = 128'h0;
  assign io_mem_acquire_bits_union = T1;
  assign T1 = 17'h1c1;
  assign io_mem_acquire_bits_a_type = T2;
  assign T2 = 3'h1;
  assign io_mem_acquire_bits_is_builtin_type = T3;
  assign T3 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T4;
  assign T4 = 2'h0;
  assign io_mem_acquire_bits_client_xact_id = T5;
  assign T5 = 6'h0;
  assign io_mem_acquire_bits_addr_block = T6;
  assign T6 = T7;
  assign T7 = refill_addr >> 3'h6;
  assign T8 = T171 ? s1_addr : refill_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T170 & T13;
  assign T13 = s1_miss ^ 1'h1;
  assign s1_miss = out_valid & T14;
  assign T14 = s1_any_tag_hit ^ 1'h1;
  assign s1_any_tag_hit = T15;
  assign T15 = T20 & T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = T18 | s1_disparity_3;
  assign s1_disparity_3 = 1'h0;
  assign T18 = T19 | s1_disparity_2;
  assign s1_disparity_2 = 1'h0;
  assign T19 = s1_disparity_0 | s1_disparity_1;
  assign s1_disparity_1 = 1'h0;
  assign s1_disparity_0 = 1'h0;
  assign T20 = T138 | s1_tag_hit_3;
  assign s1_tag_hit_3 = T21;
  assign T21 = T83 & s1_tag_match_3;
  assign s1_tag_match_3 = T22;
  assign T22 = T23 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hc];
  assign T23 = T24[7'h4f:6'h3c];
  assign T80 = T82 & s0_valid;
  assign s0_valid = io_req_valid | T81;
  assign T81 = s1_valid & stall;
  assign stall = io_resp_ready ^ 1'h1;
  assign T230 = reset ? 1'h0 : T75;
  assign T75 = T79 | T76;
  assign T76 = T78 & T77;
  assign T77 = io_req_bits_kill ^ 1'h1;
  assign T78 = s1_valid & stall;
  assign T79 = io_req_valid & rdy;
  assign T82 = refill_done ^ 1'h1;
  assign refill_done = T58 & refill_wrap;
  assign refill_wrap = T57 & T54;
  assign T54 = refill_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T55;
  assign T55 = T57 ? T56 : refill_cnt;
  assign T56 = refill_cnt + 2'h1;
  assign T57 = 1'h1 & FlowThroughSerializer_io_out_valid;
  assign T58 = state == 2'h3;
  assign T232 = reset ? 2'h0 : T59;
  assign T59 = T69 ? 2'h0 : T60;
  assign T60 = T67 ? 2'h3 : T61;
  assign T61 = T65 ? 2'h2 : T62;
  assign T62 = T63 ? 2'h1 : state;
  assign T63 = T64 & s1_miss;
  assign T64 = 2'h0 == state;
  assign T65 = T66 & io_mem_acquire_ready;
  assign T66 = 2'h1 == state;
  assign T67 = T68 & io_mem_grant_valid;
  assign T68 = 2'h2 == state;
  assign T69 = T70 & refill_done;
  assign T70 = 2'h3 == state;
  assign T73 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T74 ? s1_pgoff : io_req_bits_idx;
  assign T74 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .init(init),
    .RW0A(refill_done ? s1_idx : T73),
    .RW0E(T80 || refill_done),
    .RW0W(refill_done),
    .RW0I(T49),
    .RW0M(T26),
    .RW0O(T24)
  );
  assign T26 = T27;
  assign T27 = {T44, T28};
  assign T28 = {T42, T29};
  assign T29 = 20'h0 - T233;
  assign T233 = {19'h0, T30};
  assign T30 = repl_way == 2'h0;
  assign repl_way = R31[1'h1:1'h0];
  assign T234 = reset ? 16'h1 : T32;
  assign T32 = s1_miss ? T33 : R31;
  assign T33 = {T35, T34};
  assign T34 = R31[4'hf:1'h1];
  assign T35 = T37 ^ T36;
  assign T36 = R31[3'h5];
  assign T37 = T39 ^ T38;
  assign T38 = R31[2'h3];
  assign T39 = T41 ^ T40;
  assign T40 = R31[2'h2];
  assign T41 = R31[1'h0];
  assign T42 = 20'h0 - T235;
  assign T235 = {19'h0, T43};
  assign T43 = repl_way == 2'h1;
  assign T44 = {T47, T45};
  assign T45 = 20'h0 - T236;
  assign T236 = {19'h0, T46};
  assign T46 = repl_way == 2'h2;
  assign T47 = 20'h0 - T237;
  assign T237 = {19'h0, T48};
  assign T48 = repl_way == 2'h3;
  assign T49 = T50;
  assign T50 = {T53, T51};
  assign T51 = {T52, T52};
  assign T52 = refill_tag;
  assign refill_tag = refill_addr[5'h1f:4'hc];
  assign T53 = {T52, T52};
  assign s1_idx = s1_addr[4'hb:3'h6];
  assign T72 = T80 ? T73 : R71;
  assign T83 = T137 & T84;
  assign T84 = T85;
  assign T85 = vb_array[T86];
  assign T86 = {2'h3, T87};
  assign T87 = s1_pgoff[4'hb:3'h6];
  assign T238 = reset ? 256'h0 : T88;
  assign T88 = T136 ? T129 : T89;
  assign T89 = T128 ? T121 : T90;
  assign T90 = T120 ? T113 : T91;
  assign T91 = T112 ? T105 : T92;
  assign T92 = io_invalidate ? 256'h0 : T93;
  assign T93 = T101 ? T94 : vb_array;
  assign T94 = T99 | T95;
  assign T95 = T239 & T96;
  assign T96 = 1'h1 << T97;
  assign T97 = {repl_way, s1_idx};
  assign T239 = T98 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T98 = 1'h1;
  assign T99 = vb_array & T100;
  assign T100 = ~ T96;
  assign T101 = refill_done & T102;
  assign T102 = invalidated ^ 1'h1;
  assign T103 = T64 ? 1'h0 : T104;
  assign T104 = io_invalidate ? 1'h1 : invalidated;
  assign T105 = T110 | T240;
  assign T240 = {T242, T106};
  assign T106 = T241 & T107;
  assign T107 = 1'h1 << T108;
  assign T108 = {1'h0, s1_idx};
  assign T241 = T109 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T109 = 1'h0;
  assign T242 = T243 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T243 = T106[7'h7f];
  assign T110 = vb_array & T244;
  assign T244 = {128'h0, T111};
  assign T111 = ~ T107;
  assign T112 = s1_valid & s1_disparity_0;
  assign T113 = T118 | T245;
  assign T245 = {T247, T114};
  assign T114 = T246 & T115;
  assign T115 = 1'h1 << T116;
  assign T116 = {1'h1, s1_idx};
  assign T246 = T117 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T117 = 1'h0;
  assign T247 = T248 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T248 = T114[7'h7f];
  assign T118 = vb_array & T249;
  assign T249 = {128'h0, T119};
  assign T119 = ~ T115;
  assign T120 = s1_valid & s1_disparity_1;
  assign T121 = T126 | T122;
  assign T122 = T250 & T123;
  assign T123 = 1'h1 << T124;
  assign T124 = {2'h2, s1_idx};
  assign T250 = T125 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T125 = 1'h0;
  assign T126 = vb_array & T127;
  assign T127 = ~ T123;
  assign T128 = s1_valid & s1_disparity_2;
  assign T129 = T134 | T130;
  assign T130 = T251 & T131;
  assign T131 = 1'h1 << T132;
  assign T132 = {2'h3, s1_idx};
  assign T251 = T133 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T133 = 1'h0;
  assign T134 = vb_array & T135;
  assign T135 = ~ T131;
  assign T136 = s1_valid & s1_disparity_3;
  assign T137 = io_invalidate ^ 1'h1;
  assign T138 = T148 | s1_tag_hit_2;
  assign s1_tag_hit_2 = T139;
  assign T139 = T142 & s1_tag_match_2;
  assign s1_tag_match_2 = T140;
  assign T140 = T141 == s1_tag;
  assign T141 = T24[6'h3b:6'h28];
  assign T142 = T147 & T143;
  assign T143 = T144;
  assign T144 = vb_array[T145];
  assign T145 = {2'h2, T146};
  assign T146 = s1_pgoff[4'hb:3'h6];
  assign T147 = io_invalidate ^ 1'h1;
  assign T148 = s1_tag_hit_0 | s1_tag_hit_1;
  assign s1_tag_hit_1 = T149;
  assign T149 = T152 & s1_tag_match_1;
  assign s1_tag_match_1 = T150;
  assign T150 = T151 == s1_tag;
  assign T151 = T24[6'h27:5'h14];
  assign T152 = T157 & T153;
  assign T153 = T154;
  assign T154 = vb_array[T155];
  assign T155 = {1'h1, T156};
  assign T156 = s1_pgoff[4'hb:3'h6];
  assign T157 = io_invalidate ^ 1'h1;
  assign s1_tag_hit_0 = T158;
  assign T158 = T161 & s1_tag_match_0;
  assign s1_tag_match_0 = T159;
  assign T159 = T160 == s1_tag;
  assign T160 = T24[5'h13:1'h0];
  assign T161 = T166 & T162;
  assign T162 = T163;
  assign T163 = vb_array[T164];
  assign T164 = {1'h0, T165};
  assign T165 = s1_pgoff[4'hb:3'h6];
  assign T166 = io_invalidate ^ 1'h1;
  assign out_valid = T168 & T167;
  assign T167 = state == 2'h0;
  assign T168 = s1_valid & T169;
  assign T169 = io_req_bits_kill ^ 1'h1;
  assign T170 = state == 2'h0;
  assign T171 = T172 & s1_miss;
  assign T172 = s1_valid & T173;
  assign T173 = state == 2'h0;
  assign io_mem_acquire_valid = T174;
  assign T174 = state == 2'h1;
  assign io_resp_bits_datablock = T175;
  assign T175 = T189 | T176;
  assign T176 = s1_tag_hit_3 ? s1_dout_3 : 128'h0;
  assign s1_dout_3 = T177;
  assign T187 = T188 & s0_valid;
  assign T188 = T181 ^ 1'h1;
  assign T181 = FlowThroughSerializer_io_out_valid & T182;
  assign T182 = repl_way == 2'h3;
  assign T186 = s0_pgoff[4'hb:3'h4];
  ICache_T178 T178 (
    .CLK(clk),
    .init(init),
    .RW0A(T181 ? T183 : T186),
    .RW0E(T187 || T181),
    .RW0W(T181),
    .RW0I(T180),
    .RW0O(T177)
  );
  assign T180 = FlowThroughSerializer_io_out_bits_data;
  assign T183 = {s1_idx, refill_cnt};
  assign T185 = T187 ? T186 : R184;
  assign T189 = T203 | T190;
  assign T190 = s1_tag_hit_2 ? s1_dout_2 : 128'h0;
  assign s1_dout_2 = T191;
  assign T201 = T202 & s0_valid;
  assign T202 = T195 ^ 1'h1;
  assign T195 = FlowThroughSerializer_io_out_valid & T196;
  assign T196 = repl_way == 2'h2;
  assign T200 = s0_pgoff[4'hb:3'h4];
  ICache_T178 T192 (
    .CLK(clk),
    .init(init),
    .RW0A(T195 ? T197 : T200),
    .RW0E(T201 || T195),
    .RW0W(T195),
    .RW0I(T194),
    .RW0O(T191)
  );
  assign T194 = FlowThroughSerializer_io_out_bits_data;
  assign T197 = {s1_idx, refill_cnt};
  assign T199 = T201 ? T200 : R198;
  assign T203 = T217 | T204;
  assign T204 = s1_tag_hit_1 ? s1_dout_1 : 128'h0;
  assign s1_dout_1 = T205;
  assign T215 = T216 & s0_valid;
  assign T216 = T209 ^ 1'h1;
  assign T209 = FlowThroughSerializer_io_out_valid & T210;
  assign T210 = repl_way == 2'h1;
  assign T214 = s0_pgoff[4'hb:3'h4];
  ICache_T178 T206 (
    .CLK(clk),
    .init(init),
    .RW0A(T209 ? T211 : T214),
    .RW0E(T215 || T209),
    .RW0W(T209),
    .RW0I(T208),
    .RW0O(T205)
  );
  assign T208 = FlowThroughSerializer_io_out_bits_data;
  assign T211 = {s1_idx, refill_cnt};
  assign T213 = T215 ? T214 : R212;
  assign T217 = s1_tag_hit_0 ? s1_dout_0 : 128'h0;
  assign s1_dout_0 = T218;
  assign T228 = T229 & s0_valid;
  assign T229 = T222 ^ 1'h1;
  assign T222 = FlowThroughSerializer_io_out_valid & T223;
  assign T223 = repl_way == 2'h0;
  assign T227 = s0_pgoff[4'hb:3'h4];
  ICache_T178 T219 (
    .CLK(clk),
    .init(init),
    .RW0A(T222 ? T224 : T227),
    .RW0E(T228 || T222),
    .RW0W(T222),
    .RW0I(T221),
    .RW0O(T218)
  );
  assign T221 = FlowThroughSerializer_io_out_bits_data;
  assign T224 = {s1_idx, refill_cnt};
  assign T226 = T228 ? T227 : R225;
  assign io_resp_valid = s1_hit;
  assign s1_hit = out_valid & s1_any_tag_hit;
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       //.io_out_bits_client_xact_id(  )
       //.io_out_bits_manager_xact_id(  )
       //.io_out_bits_is_builtin_type(  )
       //.io_out_bits_g_type(  )
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );

  always @(posedge clk) begin
    if(T171) begin
      refill_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T75;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T57) begin
      refill_cnt <= T56;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T69) begin
      state <= 2'h0;
    end else if(T67) begin
      state <= 2'h3;
    end else if(T65) begin
      state <= 2'h2;
    end else if(T63) begin
      state <= 2'h1;
    end
    if(reset) begin
      R31 <= 16'h1;
    end else if(s1_miss) begin
      R31 <= T33;
    end
    if(T80) begin
      R71 <= T73;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else if(T136) begin
      vb_array <= T129;
    end else if(T128) begin
      vb_array <= T121;
    end else if(T120) begin
      vb_array <= T113;
    end else if(T112) begin
      vb_array <= T105;
    end else if(io_invalidate) begin
      vb_array <= 256'h0;
    end else if(T101) begin
      vb_array <= T94;
    end
    if(T64) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(T187) begin
      R184 <= T186;
    end
    if(T201) begin
      R198 <= T200;
    end
    if(T215) begin
      R212 <= T214;
    end
    if(T228) begin
      R225 <= T227;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input [7:0] io_clear_mask,
    input [33:0] io_tag,
    output io_hit,
    output[7:0] io_hits,
    output[7:0] io_valid_bits,
    input  io_write,
    input [33:0] io_write_tag,
    input [2:0] io_write_addr
);

  reg [7:0] vb_array;
  wire[7:0] T44;
  wire[7:0] T0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[7:0] T4;
  wire[7:0] T45;
  wire T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire[7:0] T11;
  wire[3:0] T12;
  wire[1:0] T13;
  wire hits_0;
  wire T14;
  wire[33:0] T15;
  reg [33:0] cam_tags [7:0];
  wire[33:0] T16;
  wire T17;
  wire hits_1;
  wire T18;
  wire[33:0] T19;
  wire T20;
  wire[1:0] T21;
  wire hits_2;
  wire T22;
  wire[33:0] T23;
  wire T24;
  wire hits_3;
  wire T25;
  wire[33:0] T26;
  wire T27;
  wire[3:0] T28;
  wire[1:0] T29;
  wire hits_4;
  wire T30;
  wire[33:0] T31;
  wire T32;
  wire hits_5;
  wire T33;
  wire[33:0] T34;
  wire T35;
  wire[1:0] T36;
  wire hits_6;
  wire T37;
  wire[33:0] T38;
  wire T39;
  wire hits_7;
  wire T40;
  wire[33:0] T41;
  wire T42;
  wire T43;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_valid_bits = vb_array;
  assign T44 = reset ? 8'h0 : T0;
  assign T0 = io_clear ? T8 : T1;
  assign T1 = io_write ? T2 : vb_array;
  assign T2 = T6 | T3;
  assign T3 = T45 & T4;
  assign T4 = 1'h1 << io_write_addr;
  assign T45 = T5 ? 8'hff : 8'h0;
  assign T5 = 1'h1;
  assign T6 = vb_array & T7;
  assign T7 = ~ T4;
  assign T8 = vb_array & T9;
  assign T9 = ~ io_clear_mask;
  assign io_hits = T10;
  assign T10 = T11;
  assign T11 = {T28, T12};
  assign T12 = {T21, T13};
  assign T13 = {hits_1, hits_0};
  assign hits_0 = T17 & T14;
  assign T14 = T15 == io_tag;
  assign T15 = cam_tags[3'h0];
  assign T17 = vb_array[1'h0];
  assign hits_1 = T20 & T18;
  assign T18 = T19 == io_tag;
  assign T19 = cam_tags[3'h1];
  assign T20 = vb_array[1'h1];
  assign T21 = {hits_3, hits_2};
  assign hits_2 = T24 & T22;
  assign T22 = T23 == io_tag;
  assign T23 = cam_tags[3'h2];
  assign T24 = vb_array[2'h2];
  assign hits_3 = T27 & T25;
  assign T25 = T26 == io_tag;
  assign T26 = cam_tags[3'h3];
  assign T27 = vb_array[2'h3];
  assign T28 = {T36, T29};
  assign T29 = {hits_5, hits_4};
  assign hits_4 = T32 & T30;
  assign T30 = T31 == io_tag;
  assign T31 = cam_tags[3'h4];
  assign T32 = vb_array[3'h4];
  assign hits_5 = T35 & T33;
  assign T33 = T34 == io_tag;
  assign T34 = cam_tags[3'h5];
  assign T35 = vb_array[3'h5];
  assign T36 = {hits_7, hits_6};
  assign hits_6 = T39 & T37;
  assign T37 = T38 == io_tag;
  assign T38 = cam_tags[3'h6];
  assign T39 = vb_array[3'h6];
  assign hits_7 = T42 & T40;
  assign T40 = T41 == io_tag;
  assign T41 = cam_tags[3'h7];
  assign T42 = vb_array[3'h7];
  assign io_hit = T43;
  assign T43 = io_hits != 8'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 8'h0;
    end else if(io_clear) begin
      vb_array <= T8;
    end else if(io_write) begin
      vb_array <= T2;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [27:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    input  io_req_bits_store,
    output io_resp_miss,
    output[19:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    output[7:0] io_resp_hit_idx,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate
);

  reg [2:0] r_refill_waddr;
  wire[2:0] T0;
  wire[2:0] repl_waddr;
  wire[2:0] T1;
  wire[3:0] T2;
  wire T3;
  reg [7:0] R4;
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[14:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[2:0] T479;
  wire[1:0] T480;
  wire T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[3:0] T484;
  wire[3:0] T485;
  wire[3:0] T486;
  wire[1:0] T487;
  wire T488;
  wire T489;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[7:0] T16;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[10:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[7:0] T26;
  wire T27;
  wire tlb_hit;
  wire tag_hit;
  wire[7:0] tag_hits;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] w_array;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[3:0] T33;
  wire[1:0] T34;
  reg  uw_array_0;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[7:0] T46;
  wire[2:0] T47;
  reg  uw_array_1;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  reg  uw_array_2;
  wire T52;
  wire T53;
  wire T54;
  reg  uw_array_3;
  wire T55;
  wire T56;
  wire T57;
  wire[3:0] T58;
  wire[1:0] T59;
  reg  uw_array_4;
  wire T60;
  wire T61;
  wire T62;
  reg  uw_array_5;
  wire T63;
  wire T64;
  wire T65;
  wire[1:0] T66;
  reg  uw_array_6;
  wire T67;
  wire T68;
  wire T69;
  reg  uw_array_7;
  wire T70;
  wire T71;
  wire T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire[3:0] T75;
  wire[1:0] T76;
  reg  sw_array_0;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire[2:0] T87;
  reg  sw_array_1;
  wire T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  reg  sw_array_2;
  wire T92;
  wire T93;
  wire T94;
  reg  sw_array_3;
  wire T95;
  wire T96;
  wire T97;
  wire[3:0] T98;
  wire[1:0] T99;
  reg  sw_array_4;
  wire T100;
  wire T101;
  wire T102;
  reg  sw_array_5;
  wire T103;
  wire T104;
  wire T105;
  wire[1:0] T106;
  reg  sw_array_6;
  wire T107;
  wire T108;
  wire T109;
  reg  sw_array_7;
  wire T110;
  wire T111;
  wire T112;
  wire priv_s;
  wire[1:0] priv;
  wire T113;
  wire T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[3:0] T117;
  wire[1:0] T118;
  reg  dirty_array_0;
  wire T119;
  wire T120;
  wire T121;
  wire[7:0] T122;
  wire[2:0] T123;
  reg  dirty_array_1;
  wire T124;
  wire T125;
  wire T126;
  wire[1:0] T127;
  reg  dirty_array_2;
  wire T128;
  wire T129;
  wire T130;
  reg  dirty_array_3;
  wire T131;
  wire T132;
  wire T133;
  wire[3:0] T134;
  wire[1:0] T135;
  reg  dirty_array_4;
  wire T136;
  wire T137;
  wire T138;
  reg  dirty_array_5;
  wire T139;
  wire T140;
  wire T141;
  wire[1:0] T142;
  reg  dirty_array_6;
  wire T143;
  wire T144;
  wire T145;
  reg  dirty_array_7;
  wire T146;
  wire T147;
  wire T148;
  wire vm_enabled;
  wire T149;
  wire T150;
  wire priv_uses_vm;
  wire T151;
  wire[2:0] T152;
  wire T153;
  wire[1:0] T154;
  wire T155;
  wire[2:0] T490;
  wire[2:0] T491;
  wire[2:0] T492;
  wire[2:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire[2:0] T496;
  wire T497;
  wire[7:0] T156;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire has_invalid_entry;
  wire T157;
  wire T158;
  wire tlb_miss;
  wire T159;
  wire bad_va;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[33:0] T504;
  reg [34:0] r_refill_tag;
  wire[34:0] T165;
  wire[34:0] lookup_tag;
  wire[34:0] T166;
  wire T167;
  wire T168;
  reg [1:0] state;
  wire[1:0] T505;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[33:0] T506;
  wire[7:0] T181;
  wire[7:0] T182;
  wire[7:0] T183;
  wire[7:0] T184;
  wire[7:0] T185;
  wire[7:0] T186;
  wire[7:0] T187;
  wire[3:0] T188;
  wire[1:0] T189;
  reg  valid_array_0;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[7:0] T194;
  wire[2:0] T195;
  reg  valid_array_1;
  wire T196;
  wire T197;
  wire T198;
  wire[1:0] T199;
  reg  valid_array_2;
  wire T200;
  wire T201;
  wire T202;
  reg  valid_array_3;
  wire T203;
  wire T204;
  wire T205;
  wire[3:0] T206;
  wire[1:0] T207;
  reg  valid_array_4;
  wire T208;
  wire T209;
  wire T210;
  reg  valid_array_5;
  wire T211;
  wire T212;
  wire T213;
  wire[1:0] T214;
  reg  valid_array_6;
  wire T215;
  wire T216;
  wire T217;
  reg  valid_array_7;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  reg  r_req_instruction;
  wire T223;
  reg  r_req_store;
  wire T224;
  wire[26:0] T507;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire[7:0] T230;
  wire[7:0] x_array;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[3:0] T233;
  wire[1:0] T234;
  reg  ux_array_0;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire[7:0] T246;
  wire[2:0] T247;
  reg  ux_array_1;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  reg  ux_array_2;
  wire T252;
  wire T253;
  wire T254;
  reg  ux_array_3;
  wire T255;
  wire T256;
  wire T257;
  wire[3:0] T258;
  wire[1:0] T259;
  reg  ux_array_4;
  wire T260;
  wire T261;
  wire T262;
  reg  ux_array_5;
  wire T263;
  wire T264;
  wire T265;
  wire[1:0] T266;
  reg  ux_array_6;
  wire T267;
  wire T268;
  wire T269;
  reg  ux_array_7;
  wire T270;
  wire T271;
  wire T272;
  wire[7:0] T273;
  wire[7:0] T274;
  wire[3:0] T275;
  wire[1:0] T276;
  reg  sx_array_0;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire[7:0] T286;
  wire[2:0] T287;
  reg  sx_array_1;
  wire T288;
  wire T289;
  wire T290;
  wire[1:0] T291;
  reg  sx_array_2;
  wire T292;
  wire T293;
  wire T294;
  reg  sx_array_3;
  wire T295;
  wire T296;
  wire T297;
  wire[3:0] T298;
  wire[1:0] T299;
  reg  sx_array_4;
  wire T300;
  wire T301;
  wire T302;
  reg  sx_array_5;
  wire T303;
  wire T304;
  wire T305;
  wire[1:0] T306;
  reg  sx_array_6;
  wire T307;
  wire T308;
  wire T309;
  reg  sx_array_7;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire[2:0] T317;
  wire[2:0] T318;
  wire[2:0] T319;
  wire T320;
  wire T321;
  wire[31:0] paddr;
  wire T322;
  wire[2:0] T323;
  wire[2:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire[2:0] T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire addr_ok;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire[7:0] T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire[7:0] T360;
  wire[7:0] r_array;
  wire[7:0] T361;
  wire[7:0] T362;
  wire[3:0] T363;
  wire[1:0] T364;
  reg  ur_array_0;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire[7:0] T374;
  wire[2:0] T375;
  reg  ur_array_1;
  wire T376;
  wire T377;
  wire T378;
  wire[1:0] T379;
  reg  ur_array_2;
  wire T380;
  wire T381;
  wire T382;
  reg  ur_array_3;
  wire T383;
  wire T384;
  wire T385;
  wire[3:0] T386;
  wire[1:0] T387;
  reg  ur_array_4;
  wire T388;
  wire T389;
  wire T390;
  reg  ur_array_5;
  wire T391;
  wire T392;
  wire T393;
  wire[1:0] T394;
  reg  ur_array_6;
  wire T395;
  wire T396;
  wire T397;
  reg  ur_array_7;
  wire T398;
  wire T399;
  wire T400;
  wire[7:0] T401;
  wire[7:0] T402;
  wire[3:0] T403;
  wire[1:0] T404;
  reg  sr_array_0;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[7:0] T412;
  wire[2:0] T413;
  reg  sr_array_1;
  wire T414;
  wire T415;
  wire T416;
  wire[1:0] T417;
  reg  sr_array_2;
  wire T418;
  wire T419;
  wire T420;
  reg  sr_array_3;
  wire T421;
  wire T422;
  wire T423;
  wire[3:0] T424;
  wire[1:0] T425;
  reg  sr_array_4;
  wire T426;
  wire T427;
  wire T428;
  reg  sr_array_5;
  wire T429;
  wire T430;
  wire T431;
  wire[1:0] T432;
  reg  sr_array_6;
  wire T433;
  wire T434;
  wire T435;
  reg  sr_array_7;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[19:0] T444;
  wire[19:0] T445;
  wire[19:0] T446;
  wire[19:0] T447;
  wire[19:0] T448;
  reg [19:0] tag_ram [7:0];
  wire[19:0] T449;
  wire T450;
  wire[19:0] T451;
  wire[19:0] T452;
  wire[19:0] T453;
  wire T454;
  wire[19:0] T455;
  wire[19:0] T456;
  wire[19:0] T457;
  wire T458;
  wire[19:0] T459;
  wire[19:0] T460;
  wire[19:0] T461;
  wire T462;
  wire[19:0] T463;
  wire[19:0] T464;
  wire[19:0] T465;
  wire T466;
  wire[19:0] T467;
  wire[19:0] T468;
  wire[19:0] T469;
  wire T470;
  wire[19:0] T471;
  wire[19:0] T472;
  wire[19:0] T473;
  wire T474;
  wire[19:0] T475;
  wire[19:0] T476;
  wire T477;
  wire T478;
  wire[7:0] tag_cam_io_hits;
  wire[7:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R4 = {1{$random}};
    uw_array_0 = {1{$random}};
    uw_array_1 = {1{$random}};
    uw_array_2 = {1{$random}};
    uw_array_3 = {1{$random}};
    uw_array_4 = {1{$random}};
    uw_array_5 = {1{$random}};
    uw_array_6 = {1{$random}};
    uw_array_7 = {1{$random}};
    sw_array_0 = {1{$random}};
    sw_array_1 = {1{$random}};
    sw_array_2 = {1{$random}};
    sw_array_3 = {1{$random}};
    sw_array_4 = {1{$random}};
    sw_array_5 = {1{$random}};
    sw_array_6 = {1{$random}};
    sw_array_7 = {1{$random}};
    dirty_array_0 = {1{$random}};
    dirty_array_1 = {1{$random}};
    dirty_array_2 = {1{$random}};
    dirty_array_3 = {1{$random}};
    dirty_array_4 = {1{$random}};
    dirty_array_5 = {1{$random}};
    dirty_array_6 = {1{$random}};
    dirty_array_7 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    valid_array_0 = {1{$random}};
    valid_array_1 = {1{$random}};
    valid_array_2 = {1{$random}};
    valid_array_3 = {1{$random}};
    valid_array_4 = {1{$random}};
    valid_array_5 = {1{$random}};
    valid_array_6 = {1{$random}};
    valid_array_7 = {1{$random}};
    r_req_instruction = {1{$random}};
    r_req_store = {1{$random}};
    ux_array_0 = {1{$random}};
    ux_array_1 = {1{$random}};
    ux_array_2 = {1{$random}};
    ux_array_3 = {1{$random}};
    ux_array_4 = {1{$random}};
    ux_array_5 = {1{$random}};
    ux_array_6 = {1{$random}};
    ux_array_7 = {1{$random}};
    sx_array_0 = {1{$random}};
    sx_array_1 = {1{$random}};
    sx_array_2 = {1{$random}};
    sx_array_3 = {1{$random}};
    sx_array_4 = {1{$random}};
    sx_array_5 = {1{$random}};
    sx_array_6 = {1{$random}};
    sx_array_7 = {1{$random}};
    ur_array_0 = {1{$random}};
    ur_array_1 = {1{$random}};
    ur_array_2 = {1{$random}};
    ur_array_3 = {1{$random}};
    ur_array_4 = {1{$random}};
    ur_array_5 = {1{$random}};
    ur_array_6 = {1{$random}};
    ur_array_7 = {1{$random}};
    sr_array_0 = {1{$random}};
    sr_array_1 = {1{$random}};
    sr_array_2 = {1{$random}};
    sr_array_3 = {1{$random}};
    sr_array_4 = {1{$random}};
    sr_array_5 = {1{$random}};
    sr_array_6 = {1{$random}};
    sr_array_7 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T158 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T490 : T1;
  assign T1 = T2[2'h2:1'h0];
  assign T2 = {T152, T3};
  assign T3 = R4[T152];
  assign T5 = T27 ? T6 : R4;
  assign T6 = T16 | T7;
  assign T7 = T15 ? 8'h0 : T8;
  assign T8 = T9[3'h7:1'h0];
  assign T9 = 8'h1 << T10;
  assign T10 = {T13, T11};
  assign T11 = T479[1'h1];
  assign T479 = {T489, T480};
  assign T480 = {T488, T481};
  assign T481 = T482[1'h1];
  assign T482 = T487 | T483;
  assign T483 = T484[1'h1:1'h0];
  assign T484 = T486 | T485;
  assign T485 = tag_cam_io_hits[2'h3:1'h0];
  assign T486 = tag_cam_io_hits[3'h7:3'h4];
  assign T487 = T484[2'h3:2'h2];
  assign T488 = T487 != 2'h0;
  assign T489 = T486 != 4'h0;
  assign T13 = {1'h1, T14};
  assign T14 = T479[2'h2];
  assign T15 = T479[1'h0];
  assign T16 = T18 & T17;
  assign T17 = ~ T8;
  assign T18 = T22 | T19;
  assign T19 = T11 ? 8'h0 : T20;
  assign T20 = T21[3'h7:1'h0];
  assign T21 = 8'h1 << T13;
  assign T22 = T24 & T23;
  assign T23 = ~ T20;
  assign T24 = T26 | T25;
  assign T25 = T14 ? 8'h0 : 8'h2;
  assign T26 = R4 & 8'hfd;
  assign T27 = io_req_valid & tlb_hit;
  assign tlb_hit = vm_enabled & tag_hit;
  assign tag_hit = tag_hits != 8'h0;
  assign tag_hits = tag_cam_io_hits & T28;
  assign T28 = T115 | T29;
  assign T29 = ~ T30;
  assign T30 = io_req_bits_store ? w_array : 8'h0;
  assign w_array = priv_s ? T73 : T31;
  assign T31 = T32;
  assign T32 = {T58, T33};
  assign T33 = {T51, T34};
  assign T34 = {uw_array_1, uw_array_0};
  assign T35 = T44 ? T36 : uw_array_0;
  assign T36 = T38 & T37;
  assign T37 = io_ptw_resp_bits_error ^ 1'h1;
  assign T38 = T40 & T39;
  assign T39 = io_ptw_resp_bits_pte_typ[1'h0];
  assign T40 = T42 & T41;
  assign T41 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T42 = io_ptw_resp_bits_pte_v & T43;
  assign T43 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T44 = io_ptw_resp_valid & T45;
  assign T45 = T46[1'h0];
  assign T46 = 1'h1 << T47;
  assign T47 = r_refill_waddr;
  assign T48 = T49 ? T36 : uw_array_1;
  assign T49 = io_ptw_resp_valid & T50;
  assign T50 = T46[1'h1];
  assign T51 = {uw_array_3, uw_array_2};
  assign T52 = T53 ? T36 : uw_array_2;
  assign T53 = io_ptw_resp_valid & T54;
  assign T54 = T46[2'h2];
  assign T55 = T56 ? T36 : uw_array_3;
  assign T56 = io_ptw_resp_valid & T57;
  assign T57 = T46[2'h3];
  assign T58 = {T66, T59};
  assign T59 = {uw_array_5, uw_array_4};
  assign T60 = T61 ? T36 : uw_array_4;
  assign T61 = io_ptw_resp_valid & T62;
  assign T62 = T46[3'h4];
  assign T63 = T64 ? T36 : uw_array_5;
  assign T64 = io_ptw_resp_valid & T65;
  assign T65 = T46[3'h5];
  assign T66 = {uw_array_7, uw_array_6};
  assign T67 = T68 ? T36 : uw_array_6;
  assign T68 = io_ptw_resp_valid & T69;
  assign T69 = T46[3'h6];
  assign T70 = T71 ? T36 : uw_array_7;
  assign T71 = io_ptw_resp_valid & T72;
  assign T72 = T46[3'h7];
  assign T73 = T74;
  assign T74 = {T98, T75};
  assign T75 = {T91, T76};
  assign T76 = {sw_array_1, sw_array_0};
  assign T77 = T84 ? T78 : sw_array_0;
  assign T78 = T80 & T79;
  assign T79 = io_ptw_resp_bits_error ^ 1'h1;
  assign T80 = T82 & T81;
  assign T81 = io_ptw_resp_bits_pte_typ[1'h0];
  assign T82 = io_ptw_resp_bits_pte_v & T83;
  assign T83 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T84 = io_ptw_resp_valid & T85;
  assign T85 = T86[1'h0];
  assign T86 = 1'h1 << T87;
  assign T87 = r_refill_waddr;
  assign T88 = T89 ? T78 : sw_array_1;
  assign T89 = io_ptw_resp_valid & T90;
  assign T90 = T86[1'h1];
  assign T91 = {sw_array_3, sw_array_2};
  assign T92 = T93 ? T78 : sw_array_2;
  assign T93 = io_ptw_resp_valid & T94;
  assign T94 = T86[2'h2];
  assign T95 = T96 ? T78 : sw_array_3;
  assign T96 = io_ptw_resp_valid & T97;
  assign T97 = T86[2'h3];
  assign T98 = {T106, T99};
  assign T99 = {sw_array_5, sw_array_4};
  assign T100 = T101 ? T78 : sw_array_4;
  assign T101 = io_ptw_resp_valid & T102;
  assign T102 = T86[3'h4];
  assign T103 = T104 ? T78 : sw_array_5;
  assign T104 = io_ptw_resp_valid & T105;
  assign T105 = T86[3'h5];
  assign T106 = {sw_array_7, sw_array_6};
  assign T107 = T108 ? T78 : sw_array_6;
  assign T108 = io_ptw_resp_valid & T109;
  assign T109 = T86[3'h6];
  assign T110 = T111 ? T78 : sw_array_7;
  assign T111 = io_ptw_resp_valid & T112;
  assign T112 = T86[3'h7];
  assign priv_s = priv == 2'h1;
  assign priv = T113 ? io_ptw_status_prv1 : io_ptw_status_prv;
  assign T113 = io_ptw_status_mprv & T114;
  assign T114 = io_req_bits_instruction ^ 1'h1;
  assign T115 = T116;
  assign T116 = {T134, T117};
  assign T117 = {T127, T118};
  assign T118 = {dirty_array_1, dirty_array_0};
  assign T119 = T120 ? io_ptw_resp_bits_pte_d : dirty_array_0;
  assign T120 = io_ptw_resp_valid & T121;
  assign T121 = T122[1'h0];
  assign T122 = 1'h1 << T123;
  assign T123 = r_refill_waddr;
  assign T124 = T125 ? io_ptw_resp_bits_pte_d : dirty_array_1;
  assign T125 = io_ptw_resp_valid & T126;
  assign T126 = T122[1'h1];
  assign T127 = {dirty_array_3, dirty_array_2};
  assign T128 = T129 ? io_ptw_resp_bits_pte_d : dirty_array_2;
  assign T129 = io_ptw_resp_valid & T130;
  assign T130 = T122[2'h2];
  assign T131 = T132 ? io_ptw_resp_bits_pte_d : dirty_array_3;
  assign T132 = io_ptw_resp_valid & T133;
  assign T133 = T122[2'h3];
  assign T134 = {T142, T135};
  assign T135 = {dirty_array_5, dirty_array_4};
  assign T136 = T137 ? io_ptw_resp_bits_pte_d : dirty_array_4;
  assign T137 = io_ptw_resp_valid & T138;
  assign T138 = T122[3'h4];
  assign T139 = T140 ? io_ptw_resp_bits_pte_d : dirty_array_5;
  assign T140 = io_ptw_resp_valid & T141;
  assign T141 = T122[3'h5];
  assign T142 = {dirty_array_7, dirty_array_6};
  assign T143 = T144 ? io_ptw_resp_bits_pte_d : dirty_array_6;
  assign T144 = io_ptw_resp_valid & T145;
  assign T145 = T122[3'h6];
  assign T146 = T147 ? io_ptw_resp_bits_pte_d : dirty_array_7;
  assign T147 = io_ptw_resp_valid & T148;
  assign T148 = T122[3'h7];
  assign vm_enabled = T150 & T149;
  assign T149 = io_req_bits_passthrough ^ 1'h1;
  assign T150 = T151 & priv_uses_vm;
  assign priv_uses_vm = priv <= 2'h1;
  assign T151 = io_ptw_status_vm[2'h3];
  assign T152 = {T154, T153};
  assign T153 = R4[T154];
  assign T154 = {1'h1, T155};
  assign T155 = R4[1'h1];
  assign T490 = T503 ? 1'h0 : T491;
  assign T491 = T502 ? 1'h1 : T492;
  assign T492 = T501 ? 2'h2 : T493;
  assign T493 = T500 ? 2'h3 : T494;
  assign T494 = T499 ? 3'h4 : T495;
  assign T495 = T498 ? 3'h5 : T496;
  assign T496 = T497 ? 3'h6 : 3'h7;
  assign T497 = T156[3'h6];
  assign T156 = ~ tag_cam_io_valid_bits;
  assign T498 = T156[3'h5];
  assign T499 = T156[3'h4];
  assign T500 = T156[2'h3];
  assign T501 = T156[2'h2];
  assign T502 = T156[1'h1];
  assign T503 = T156[1'h0];
  assign has_invalid_entry = T157 ^ 1'h1;
  assign T157 = tag_cam_io_valid_bits == 8'hff;
  assign T158 = T164 & tlb_miss;
  assign tlb_miss = T162 & T159;
  assign T159 = bad_va ^ 1'h1;
  assign bad_va = T161 != T160;
  assign T160 = io_req_bits_vpn[5'h1a];
  assign T161 = io_req_bits_vpn[5'h1b];
  assign T162 = vm_enabled & T163;
  assign T163 = tag_hit ^ 1'h1;
  assign T164 = io_req_ready & io_req_valid;
  assign T504 = r_refill_tag[6'h21:1'h0];
  assign T165 = T158 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T166;
  assign T166 = {io_req_bits_asid, io_req_bits_vpn};
  assign T167 = T168 & io_ptw_resp_valid;
  assign T168 = state == 2'h2;
  assign T505 = reset ? 2'h0 : T169;
  assign T169 = io_ptw_resp_valid ? 2'h0 : T170;
  assign T170 = T179 ? 2'h3 : T171;
  assign T171 = T178 ? 2'h3 : T172;
  assign T172 = T177 ? 2'h2 : T173;
  assign T173 = T175 ? 2'h0 : T174;
  assign T174 = T158 ? 2'h1 : state;
  assign T175 = T176 & io_ptw_invalidate;
  assign T176 = state == 2'h1;
  assign T177 = T176 & io_ptw_req_ready;
  assign T178 = T177 & io_ptw_invalidate;
  assign T179 = T180 & io_ptw_invalidate;
  assign T180 = state == 2'h2;
  assign T506 = lookup_tag[6'h21:1'h0];
  assign T181 = io_ptw_invalidate ? 8'hff : T182;
  assign T182 = T185 | T183;
  assign T183 = tag_cam_io_hits & T184;
  assign T184 = ~ tag_hits;
  assign T185 = ~ T186;
  assign T186 = T187;
  assign T187 = {T206, T188};
  assign T188 = {T199, T189};
  assign T189 = {valid_array_1, valid_array_0};
  assign T190 = T192 ? T191 : valid_array_0;
  assign T191 = io_ptw_resp_bits_error ^ 1'h1;
  assign T192 = io_ptw_resp_valid & T193;
  assign T193 = T194[1'h0];
  assign T194 = 1'h1 << T195;
  assign T195 = r_refill_waddr;
  assign T196 = T197 ? T191 : valid_array_1;
  assign T197 = io_ptw_resp_valid & T198;
  assign T198 = T194[1'h1];
  assign T199 = {valid_array_3, valid_array_2};
  assign T200 = T201 ? T191 : valid_array_2;
  assign T201 = io_ptw_resp_valid & T202;
  assign T202 = T194[2'h2];
  assign T203 = T204 ? T191 : valid_array_3;
  assign T204 = io_ptw_resp_valid & T205;
  assign T205 = T194[2'h3];
  assign T206 = {T214, T207};
  assign T207 = {valid_array_5, valid_array_4};
  assign T208 = T209 ? T191 : valid_array_4;
  assign T209 = io_ptw_resp_valid & T210;
  assign T210 = T194[3'h4];
  assign T211 = T212 ? T191 : valid_array_5;
  assign T212 = io_ptw_resp_valid & T213;
  assign T213 = T194[3'h5];
  assign T214 = {valid_array_7, valid_array_6};
  assign T215 = T216 ? T191 : valid_array_6;
  assign T216 = io_ptw_resp_valid & T217;
  assign T217 = T194[3'h6];
  assign T218 = T219 ? T191 : valid_array_7;
  assign T219 = io_ptw_resp_valid & T220;
  assign T220 = T194[3'h7];
  assign T221 = io_ptw_invalidate | T222;
  assign T222 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T223 = T158 ? io_req_bits_instruction : r_req_instruction;
  assign io_ptw_req_bits_store = r_req_store;
  assign T224 = T158 ? io_req_bits_store : r_req_store;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_addr = T507;
  assign T507 = r_refill_tag[5'h1a:1'h0];
  assign io_ptw_req_valid = T225;
  assign T225 = state == 2'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_xcpt_if = T226;
  assign T226 = T313 | T227;
  assign T227 = tlb_hit & T228;
  assign T228 = T229 ^ 1'h1;
  assign T229 = T230 != 8'h0;
  assign T230 = x_array & tag_cam_io_hits;
  assign x_array = priv_s ? T273 : T231;
  assign T231 = T232;
  assign T232 = {T258, T233};
  assign T233 = {T251, T234};
  assign T234 = {ux_array_1, ux_array_0};
  assign T235 = T244 ? T236 : ux_array_0;
  assign T236 = T238 & T237;
  assign T237 = io_ptw_resp_bits_error ^ 1'h1;
  assign T238 = T240 & T239;
  assign T239 = io_ptw_resp_bits_pte_typ[1'h1];
  assign T240 = T242 & T241;
  assign T241 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T242 = io_ptw_resp_bits_pte_v & T243;
  assign T243 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T244 = io_ptw_resp_valid & T245;
  assign T245 = T246[1'h0];
  assign T246 = 1'h1 << T247;
  assign T247 = r_refill_waddr;
  assign T248 = T249 ? T236 : ux_array_1;
  assign T249 = io_ptw_resp_valid & T250;
  assign T250 = T246[1'h1];
  assign T251 = {ux_array_3, ux_array_2};
  assign T252 = T253 ? T236 : ux_array_2;
  assign T253 = io_ptw_resp_valid & T254;
  assign T254 = T246[2'h2];
  assign T255 = T256 ? T236 : ux_array_3;
  assign T256 = io_ptw_resp_valid & T257;
  assign T257 = T246[2'h3];
  assign T258 = {T266, T259};
  assign T259 = {ux_array_5, ux_array_4};
  assign T260 = T261 ? T236 : ux_array_4;
  assign T261 = io_ptw_resp_valid & T262;
  assign T262 = T246[3'h4];
  assign T263 = T264 ? T236 : ux_array_5;
  assign T264 = io_ptw_resp_valid & T265;
  assign T265 = T246[3'h5];
  assign T266 = {ux_array_7, ux_array_6};
  assign T267 = T268 ? T236 : ux_array_6;
  assign T268 = io_ptw_resp_valid & T269;
  assign T269 = T246[3'h6];
  assign T270 = T271 ? T236 : ux_array_7;
  assign T271 = io_ptw_resp_valid & T272;
  assign T272 = T246[3'h7];
  assign T273 = T274;
  assign T274 = {T298, T275};
  assign T275 = {T291, T276};
  assign T276 = {sx_array_1, sx_array_0};
  assign T277 = T284 ? T278 : sx_array_0;
  assign T278 = T280 & T279;
  assign T279 = io_ptw_resp_bits_error ^ 1'h1;
  assign T280 = T282 & T281;
  assign T281 = io_ptw_resp_bits_pte_typ[1'h1];
  assign T282 = io_ptw_resp_bits_pte_v & T283;
  assign T283 = 4'h4 <= io_ptw_resp_bits_pte_typ;
  assign T284 = io_ptw_resp_valid & T285;
  assign T285 = T286[1'h0];
  assign T286 = 1'h1 << T287;
  assign T287 = r_refill_waddr;
  assign T288 = T289 ? T278 : sx_array_1;
  assign T289 = io_ptw_resp_valid & T290;
  assign T290 = T286[1'h1];
  assign T291 = {sx_array_3, sx_array_2};
  assign T292 = T293 ? T278 : sx_array_2;
  assign T293 = io_ptw_resp_valid & T294;
  assign T294 = T286[2'h2];
  assign T295 = T296 ? T278 : sx_array_3;
  assign T296 = io_ptw_resp_valid & T297;
  assign T297 = T286[2'h3];
  assign T298 = {T306, T299};
  assign T299 = {sx_array_5, sx_array_4};
  assign T300 = T301 ? T278 : sx_array_4;
  assign T301 = io_ptw_resp_valid & T302;
  assign T302 = T286[3'h4];
  assign T303 = T304 ? T278 : sx_array_5;
  assign T304 = io_ptw_resp_valid & T305;
  assign T305 = T286[3'h5];
  assign T306 = {sx_array_7, sx_array_6};
  assign T307 = T308 ? T278 : sx_array_6;
  assign T308 = io_ptw_resp_valid & T309;
  assign T309 = T286[3'h6];
  assign T310 = T311 ? T278 : sx_array_7;
  assign T311 = io_ptw_resp_valid & T312;
  assign T312 = T286[3'h7];
  assign T313 = T314 | bad_va;
  assign T314 = T333 | T315;
  assign T315 = T316 ^ 1'h1;
  assign T316 = T317[2'h2];
  assign T317 = T332 ? 3'h7 : T318;
  assign T318 = T323 | T319;
  assign T319 = T320 ? 3'h3 : 3'h0;
  assign T320 = T322 & T321;
  assign T321 = paddr < 32'h40010200;
  assign paddr = {io_resp_ppn, 12'h0};
  assign T322 = 32'h40010000 <= paddr;
  assign T323 = T328 | T324;
  assign T324 = T325 ? 3'h3 : 3'h0;
  assign T325 = T327 & T326;
  assign T326 = paddr < 32'h40010000;
  assign T327 = 32'h40008000 <= paddr;
  assign T328 = T329 ? 3'h1 : 3'h0;
  assign T329 = T331 & T330;
  assign T330 = paddr < 32'h40008000;
  assign T331 = 32'h40000000 <= paddr;
  assign T332 = paddr < 32'h40000000;
  assign T333 = addr_ok ^ 1'h1;
  assign addr_ok = T345 | T334;
  assign T334 = T338 | T335;
  assign T335 = T337 & T336;
  assign T336 = paddr < 32'h40010200;
  assign T337 = 32'h40010000 <= paddr;
  assign T338 = T342 | T339;
  assign T339 = T341 & T340;
  assign T340 = paddr < 32'h40010000;
  assign T341 = 32'h40008000 <= paddr;
  assign T342 = T344 & T343;
  assign T343 = paddr < 32'h40008000;
  assign T344 = 32'h40000000 <= paddr;
  assign T345 = paddr < 32'h40000000;
  assign io_resp_xcpt_st = T346;
  assign T346 = T351 | T347;
  assign T347 = tlb_hit & T348;
  assign T348 = T349 ^ 1'h1;
  assign T349 = T350 != 8'h0;
  assign T350 = w_array & tag_cam_io_hits;
  assign T351 = T352 | bad_va;
  assign T352 = T355 | T353;
  assign T353 = T354 ^ 1'h1;
  assign T354 = T317[1'h1];
  assign T355 = addr_ok ^ 1'h1;
  assign io_resp_xcpt_ld = T356;
  assign T356 = T439 | T357;
  assign T357 = tlb_hit & T358;
  assign T358 = T359 ^ 1'h1;
  assign T359 = T360 != 8'h0;
  assign T360 = r_array & tag_cam_io_hits;
  assign r_array = priv_s ? T401 : T361;
  assign T361 = T362;
  assign T362 = {T386, T363};
  assign T363 = {T379, T364};
  assign T364 = {ur_array_1, ur_array_0};
  assign T365 = T372 ? T366 : ur_array_0;
  assign T366 = T368 & T367;
  assign T367 = io_ptw_resp_bits_error ^ 1'h1;
  assign T368 = T370 & T369;
  assign T369 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T370 = io_ptw_resp_bits_pte_v & T371;
  assign T371 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T372 = io_ptw_resp_valid & T373;
  assign T373 = T374[1'h0];
  assign T374 = 1'h1 << T375;
  assign T375 = r_refill_waddr;
  assign T376 = T377 ? T366 : ur_array_1;
  assign T377 = io_ptw_resp_valid & T378;
  assign T378 = T374[1'h1];
  assign T379 = {ur_array_3, ur_array_2};
  assign T380 = T381 ? T366 : ur_array_2;
  assign T381 = io_ptw_resp_valid & T382;
  assign T382 = T374[2'h2];
  assign T383 = T384 ? T366 : ur_array_3;
  assign T384 = io_ptw_resp_valid & T385;
  assign T385 = T374[2'h3];
  assign T386 = {T394, T387};
  assign T387 = {ur_array_5, ur_array_4};
  assign T388 = T389 ? T366 : ur_array_4;
  assign T389 = io_ptw_resp_valid & T390;
  assign T390 = T374[3'h4];
  assign T391 = T392 ? T366 : ur_array_5;
  assign T392 = io_ptw_resp_valid & T393;
  assign T393 = T374[3'h5];
  assign T394 = {ur_array_7, ur_array_6};
  assign T395 = T396 ? T366 : ur_array_6;
  assign T396 = io_ptw_resp_valid & T397;
  assign T397 = T374[3'h6];
  assign T398 = T399 ? T366 : ur_array_7;
  assign T399 = io_ptw_resp_valid & T400;
  assign T400 = T374[3'h7];
  assign T401 = T402;
  assign T402 = {T424, T403};
  assign T403 = {T417, T404};
  assign T404 = {sr_array_1, sr_array_0};
  assign T405 = T410 ? T406 : sr_array_0;
  assign T406 = T408 & T407;
  assign T407 = io_ptw_resp_bits_error ^ 1'h1;
  assign T408 = io_ptw_resp_bits_pte_v & T409;
  assign T409 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T410 = io_ptw_resp_valid & T411;
  assign T411 = T412[1'h0];
  assign T412 = 1'h1 << T413;
  assign T413 = r_refill_waddr;
  assign T414 = T415 ? T406 : sr_array_1;
  assign T415 = io_ptw_resp_valid & T416;
  assign T416 = T412[1'h1];
  assign T417 = {sr_array_3, sr_array_2};
  assign T418 = T419 ? T406 : sr_array_2;
  assign T419 = io_ptw_resp_valid & T420;
  assign T420 = T412[2'h2];
  assign T421 = T422 ? T406 : sr_array_3;
  assign T422 = io_ptw_resp_valid & T423;
  assign T423 = T412[2'h3];
  assign T424 = {T432, T425};
  assign T425 = {sr_array_5, sr_array_4};
  assign T426 = T427 ? T406 : sr_array_4;
  assign T427 = io_ptw_resp_valid & T428;
  assign T428 = T412[3'h4];
  assign T429 = T430 ? T406 : sr_array_5;
  assign T430 = io_ptw_resp_valid & T431;
  assign T431 = T412[3'h5];
  assign T432 = {sr_array_7, sr_array_6};
  assign T433 = T434 ? T406 : sr_array_6;
  assign T434 = io_ptw_resp_valid & T435;
  assign T435 = T412[3'h6];
  assign T436 = T437 ? T406 : sr_array_7;
  assign T437 = io_ptw_resp_valid & T438;
  assign T438 = T412[3'h7];
  assign T439 = T440 | bad_va;
  assign T440 = T443 | T441;
  assign T441 = T442 ^ 1'h1;
  assign T442 = T317[1'h0];
  assign T443 = addr_ok ^ 1'h1;
  assign io_resp_ppn = T444;
  assign T444 = vm_enabled ? T446 : T445;
  assign T445 = io_req_bits_vpn[5'h13:1'h0];
  assign T446 = T451 | T447;
  assign T447 = T450 ? T448 : 20'h0;
  assign T448 = tag_ram[3'h7];
  assign T450 = tag_cam_io_hits[3'h7];
  assign T451 = T455 | T452;
  assign T452 = T454 ? T453 : 20'h0;
  assign T453 = tag_ram[3'h6];
  assign T454 = tag_cam_io_hits[3'h6];
  assign T455 = T459 | T456;
  assign T456 = T458 ? T457 : 20'h0;
  assign T457 = tag_ram[3'h5];
  assign T458 = tag_cam_io_hits[3'h5];
  assign T459 = T463 | T460;
  assign T460 = T462 ? T461 : 20'h0;
  assign T461 = tag_ram[3'h4];
  assign T462 = tag_cam_io_hits[3'h4];
  assign T463 = T467 | T464;
  assign T464 = T466 ? T465 : 20'h0;
  assign T465 = tag_ram[3'h3];
  assign T466 = tag_cam_io_hits[2'h3];
  assign T467 = T471 | T468;
  assign T468 = T470 ? T469 : 20'h0;
  assign T469 = tag_ram[3'h2];
  assign T470 = tag_cam_io_hits[2'h2];
  assign T471 = T475 | T472;
  assign T472 = T474 ? T473 : 20'h0;
  assign T473 = tag_ram[3'h1];
  assign T474 = tag_cam_io_hits[1'h1];
  assign T475 = T477 ? T476 : 20'h0;
  assign T476 = tag_ram[3'h0];
  assign T477 = tag_cam_io_hits[1'h0];
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T478;
  assign T478 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( T221 ),
       .io_clear_mask( T181 ),
       .io_tag( T506 ),
       //.io_hit(  )
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T167 ),
       .io_write_tag( T504 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T158) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T27) begin
      R4 <= T6;
    end
    if(T44) begin
      uw_array_0 <= T36;
    end
    if(T49) begin
      uw_array_1 <= T36;
    end
    if(T53) begin
      uw_array_2 <= T36;
    end
    if(T56) begin
      uw_array_3 <= T36;
    end
    if(T61) begin
      uw_array_4 <= T36;
    end
    if(T64) begin
      uw_array_5 <= T36;
    end
    if(T68) begin
      uw_array_6 <= T36;
    end
    if(T71) begin
      uw_array_7 <= T36;
    end
    if(T84) begin
      sw_array_0 <= T78;
    end
    if(T89) begin
      sw_array_1 <= T78;
    end
    if(T93) begin
      sw_array_2 <= T78;
    end
    if(T96) begin
      sw_array_3 <= T78;
    end
    if(T101) begin
      sw_array_4 <= T78;
    end
    if(T104) begin
      sw_array_5 <= T78;
    end
    if(T108) begin
      sw_array_6 <= T78;
    end
    if(T111) begin
      sw_array_7 <= T78;
    end
    if(T120) begin
      dirty_array_0 <= io_ptw_resp_bits_pte_d;
    end
    if(T125) begin
      dirty_array_1 <= io_ptw_resp_bits_pte_d;
    end
    if(T129) begin
      dirty_array_2 <= io_ptw_resp_bits_pte_d;
    end
    if(T132) begin
      dirty_array_3 <= io_ptw_resp_bits_pte_d;
    end
    if(T137) begin
      dirty_array_4 <= io_ptw_resp_bits_pte_d;
    end
    if(T140) begin
      dirty_array_5 <= io_ptw_resp_bits_pte_d;
    end
    if(T144) begin
      dirty_array_6 <= io_ptw_resp_bits_pte_d;
    end
    if(T147) begin
      dirty_array_7 <= io_ptw_resp_bits_pte_d;
    end
    if(T158) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T179) begin
      state <= 2'h3;
    end else if(T178) begin
      state <= 2'h3;
    end else if(T177) begin
      state <= 2'h2;
    end else if(T175) begin
      state <= 2'h0;
    end else if(T158) begin
      state <= 2'h1;
    end
    if(T192) begin
      valid_array_0 <= T191;
    end
    if(T197) begin
      valid_array_1 <= T191;
    end
    if(T201) begin
      valid_array_2 <= T191;
    end
    if(T204) begin
      valid_array_3 <= T191;
    end
    if(T209) begin
      valid_array_4 <= T191;
    end
    if(T212) begin
      valid_array_5 <= T191;
    end
    if(T216) begin
      valid_array_6 <= T191;
    end
    if(T219) begin
      valid_array_7 <= T191;
    end
    if(T158) begin
      r_req_instruction <= io_req_bits_instruction;
    end
    if(T158) begin
      r_req_store <= io_req_bits_store;
    end
    if(T244) begin
      ux_array_0 <= T236;
    end
    if(T249) begin
      ux_array_1 <= T236;
    end
    if(T253) begin
      ux_array_2 <= T236;
    end
    if(T256) begin
      ux_array_3 <= T236;
    end
    if(T261) begin
      ux_array_4 <= T236;
    end
    if(T264) begin
      ux_array_5 <= T236;
    end
    if(T268) begin
      ux_array_6 <= T236;
    end
    if(T271) begin
      ux_array_7 <= T236;
    end
    if(T284) begin
      sx_array_0 <= T278;
    end
    if(T289) begin
      sx_array_1 <= T278;
    end
    if(T293) begin
      sx_array_2 <= T278;
    end
    if(T296) begin
      sx_array_3 <= T278;
    end
    if(T301) begin
      sx_array_4 <= T278;
    end
    if(T304) begin
      sx_array_5 <= T278;
    end
    if(T308) begin
      sx_array_6 <= T278;
    end
    if(T311) begin
      sx_array_7 <= T278;
    end
    if(T372) begin
      ur_array_0 <= T366;
    end
    if(T377) begin
      ur_array_1 <= T366;
    end
    if(T381) begin
      ur_array_2 <= T366;
    end
    if(T384) begin
      ur_array_3 <= T366;
    end
    if(T389) begin
      ur_array_4 <= T366;
    end
    if(T392) begin
      ur_array_5 <= T366;
    end
    if(T396) begin
      ur_array_6 <= T366;
    end
    if(T399) begin
      ur_array_7 <= T366;
    end
    if(T410) begin
      sr_array_0 <= T406;
    end
    if(T415) begin
      sr_array_1 <= T406;
    end
    if(T419) begin
      sr_array_2 <= T406;
    end
    if(T422) begin
      sr_array_3 <= T406;
    end
    if(T427) begin
      sr_array_4 <= T406;
    end
    if(T430) begin
      sr_array_5 <= T406;
    end
    if(T434) begin
      sr_array_6 <= T406;
    end
    if(T437) begin
      sr_array_7 <= T406;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_pte_ppn;
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_data,
    input [127:0] io_enq_bits_datablock,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_data,
    output[127:0] io_deq_bits_datablock,
    output io_count
);

  wire T12;
  wire[1:0] T0;
  reg  full;
  wire T13;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[159:0] T4;
  reg [159:0] ram [0:0];
  wire[159:0] T5;
  wire[159:0] T6;
  wire[159:0] T7;
  wire[31:0] T8;
  wire T9;
  wire empty;
  wire T10;
  wire T11;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T12;
  assign T12 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T13 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_datablock = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_data, io_enq_bits_datablock};
  assign io_deq_bits_data = T8;
  assign T8 = T4[8'h9f:8'h80];
  assign io_deq_valid = T9;
  assign T9 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T10;
  assign T10 = T11 | io_deq_ready;
  assign T11 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data_0,
    output io_cpu_resp_bits_mask,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output io_cpu_btb_resp_bits_mask,
    output io_cpu_btb_resp_bits_bridx,
    output[38:0] io_cpu_btb_resp_bits_target,
    output[5:0] io_cpu_btb_resp_bits_entry,
    output[6:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input  io_cpu_btb_update_bits_prediction_bits_mask,
    input  io_cpu_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_btb_update_bits_pc,
    input [38:0] io_cpu_btb_update_bits_target,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isReturn,
    input [38:0] io_cpu_btb_update_bits_br_pc,
    input  io_cpu_bht_update_valid,
    input  io_cpu_bht_update_bits_prediction_valid,
    input  io_cpu_bht_update_bits_prediction_bits_taken,
    input  io_cpu_bht_update_bits_prediction_bits_mask,
    input  io_cpu_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_bht_update_bits_prediction_bits_target,
    input [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_bht_update_bits_pc,
    input  io_cpu_bht_update_bits_taken,
    input  io_cpu_bht_update_bits_mispredict,
    input  io_cpu_ras_update_valid,
    input  io_cpu_ras_update_bits_isCall,
    input  io_cpu_ras_update_bits_isReturn,
    input [38:0] io_cpu_ras_update_bits_returnAddr,
    input  io_cpu_ras_update_bits_prediction_valid,
    input  io_cpu_ras_update_bits_prediction_bits_taken,
    input  io_cpu_ras_update_bits_prediction_bits_mask,
    input  io_cpu_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_ras_update_bits_prediction_bits_target,
    input [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
    input  io_cpu_invalidate,
    output[39:0] io_cpu_npc,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[5:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  init
);

  wire T0;
  wire T1;
  reg  s1_same_block;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire s0_same_block;
  wire T6;
  wire[39:0] T7;
  wire[39:0] s1_pc;
  wire[39:0] T8;
  wire[39:0] T9;
  reg [39:0] s1_pc_;
  wire[39:0] T10;
  wire[39:0] T11;
  wire[39:0] npc;
  wire[39:0] T12;
  wire[39:0] predicted_npc;
  wire[39:0] ntpc;
  wire[38:0] T13;
  wire[36:0] T14;
  wire[39:0] ntpc_0;
  wire T15;
  wire T16;
  wire T17;
  wire[39:0] btbTarget;
  wire T18;
  reg [39:0] s2_pc;
  wire[39:0] T68;
  wire[39:0] T19;
  wire T20;
  wire T21;
  wire icmiss;
  wire T22;
  wire s2_resp_valid;
  reg  s2_valid;
  wire T69;
  wire T23;
  wire T24;
  wire T25;
  wire[39:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire stall;
  wire T33;
  wire T34;
  wire[27:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[11:0] T70;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[38:0] T71;
  wire T47;
  wire T48;
  wire T49;
  wire[39:0] T50;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T51;
  wire T52;
  reg [6:0] s2_btb_resp_bits_bht_history;
  wire[6:0] T53;
  reg [5:0] s2_btb_resp_bits_entry;
  wire[5:0] T54;
  reg [38:0] s2_btb_resp_bits_target;
  wire[38:0] T55;
  reg  s2_btb_resp_bits_bridx;
  wire T56;
  reg  s2_btb_resp_bits_mask;
  wire T57;
  reg  s2_btb_resp_bits_taken;
  wire T58;
  reg  s2_btb_resp_valid;
  wire T72;
  wire T59;
  reg  s2_xcpt_if;
  wire T73;
  wire T60;
  wire T74;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T75;
  wire[31:0] T63;
  wire[127:0] fetch_data;
  wire[6:0] T64;
  wire[1:0] T65;
  wire[127:0] s2_resp_data;
  wire T66;
  wire T67;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire btb_io_resp_bits_mask;
  wire btb_io_resp_bits_bridx;
  wire[38:0] btb_io_resp_bits_target;
  wire[5:0] btb_io_resp_bits_entry;
  wire[6:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[127:0] Queue_io_deq_bits_datablock;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[5:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire tlb_io_resp_miss;
  wire[19:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[26:0] tlb_io_ptw_req_bits_addr;
  wire[1:0] tlb_io_ptw_req_bits_prv;
  wire tlb_io_ptw_req_bits_store;
  wire tlb_io_ptw_req_bits_fetch;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s1_same_block = {1{$random}};
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_bridx = {1{$random}};
    s2_btb_resp_bits_mask = {1{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T34 & T1;
  assign T1 = s1_same_block ^ 1'h1;
  assign T2 = io_cpu_req_valid ? 1'h0 : T3;
  assign T3 = T32 ? T4 : s1_same_block;
  assign T4 = s0_same_block & T5;
  assign T5 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T27 & T6;
  assign T6 = T26 == T7;
  assign T7 = s1_pc & 40'h10;
  assign s1_pc = ~ T8;
  assign T8 = T9 | 40'h3;
  assign T9 = ~ s1_pc_;
  assign T10 = io_cpu_req_valid ? io_cpu_req_bits_pc : T11;
  assign T11 = T32 ? npc : s1_pc_;
  assign npc = T12;
  assign T12 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : ntpc;
  assign ntpc = {T15, T13};
  assign T13 = {T14, 2'h0};
  assign T14 = ntpc_0[6'h26:2'h2];
  assign ntpc_0 = s1_pc + 40'h4;
  assign T15 = T17 & T16;
  assign T16 = ntpc_0[6'h26];
  assign T17 = s1_pc[6'h26];
  assign btbTarget = {T18, btb_io_resp_bits_target};
  assign T18 = btb_io_resp_bits_target[6'h26];
  assign T68 = reset ? 40'h200 : T19;
  assign T19 = T20 ? s1_pc : s2_pc;
  assign T20 = T32 & T21;
  assign T21 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T22;
  assign T22 = s2_resp_valid ^ 1'h1;
  assign s2_resp_valid = Queue_io_deq_valid;
  assign T69 = reset ? 1'h1 : T23;
  assign T23 = io_cpu_req_valid ? 1'h0 : T24;
  assign T24 = T32 ? T25 : s2_valid;
  assign T25 = icmiss ^ 1'h1;
  assign T26 = ntpc & 40'h10;
  assign T27 = T29 & T28;
  assign T28 = btb_io_resp_bits_taken ^ 1'h1;
  assign T29 = T31 & T30;
  assign T30 = io_cpu_req_valid ^ 1'h1;
  assign T31 = icmiss ^ 1'h1;
  assign T32 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T33;
  assign T33 = io_cpu_resp_ready ^ 1'h1;
  assign T34 = stall ^ 1'h1;
  assign T35 = s1_pc >> 4'hc;
  assign T36 = T38 & T37;
  assign T37 = icmiss ^ 1'h1;
  assign T38 = stall ^ 1'h1;
  assign T39 = T40 | io_ptw_invalidate;
  assign T40 = T41 | icmiss;
  assign T41 = T42 | tlb_io_resp_xcpt_if;
  assign T42 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T70 = io_cpu_npc[4'hb:1'h0];
  assign T43 = T45 & T44;
  assign T44 = s0_same_block ^ 1'h1;
  assign T45 = stall ^ 1'h1;
  assign T46 = io_cpu_invalidate | io_ptw_invalidate;
  assign T71 = s1_pc[6'h26:1'h0];
  assign T47 = T49 & T48;
  assign T48 = icmiss ^ 1'h1;
  assign T49 = stall ^ 1'h1;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_npc = T50;
  assign T50 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T51 = T52 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T52 = T20 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T53 = T52 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T54 = T52 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T55 = T52 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign T56 = T52 ? btb_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign T57 = T52 ? btb_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T58 = T52 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T72 = reset ? 1'h0 : T59;
  assign T59 = T20 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T73 = reset ? 1'h0 : T60;
  assign T60 = T20 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_mask = T74;
  assign T74 = T61[1'h0];
  assign T61 = s2_btb_resp_valid ? T62 : 2'h3;
  assign T62 = 2'h3 & T75;
  assign T75 = {1'h0, s2_btb_resp_bits_mask};
  assign io_cpu_resp_bits_data_0 = T63;
  assign T63 = fetch_data[5'h1f:1'h0];
  assign fetch_data = s2_resp_data >> T64;
  assign T64 = T65 << 3'h5;
  assign T65 = s2_pc[2'h3:2'h2];
  assign s2_resp_data = Queue_io_deq_bits_datablock;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_valid = T66;
  assign T66 = s2_valid & T67;
  assign T67 = s2_xcpt_if | s2_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T47 ),
       .io_req_bits_addr( T71 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_mask( btb_io_resp_bits_mask ),
       .io_resp_bits_bridx( btb_io_resp_bits_bridx ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_btb_update_valid( io_cpu_btb_update_valid ),
       .io_btb_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_btb_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_btb_update_bits_prediction_bits_mask( io_cpu_btb_update_bits_prediction_bits_mask ),
       .io_btb_update_bits_prediction_bits_bridx( io_cpu_btb_update_bits_prediction_bits_bridx ),
       .io_btb_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_btb_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_btb_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_btb_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_btb_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_btb_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_btb_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_btb_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_btb_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_btb_update_bits_br_pc( io_cpu_btb_update_bits_br_pc ),
       .io_bht_update_valid( io_cpu_bht_update_valid ),
       .io_bht_update_bits_prediction_valid( io_cpu_bht_update_bits_prediction_valid ),
       .io_bht_update_bits_prediction_bits_taken( io_cpu_bht_update_bits_prediction_bits_taken ),
       .io_bht_update_bits_prediction_bits_mask( io_cpu_bht_update_bits_prediction_bits_mask ),
       .io_bht_update_bits_prediction_bits_bridx( io_cpu_bht_update_bits_prediction_bits_bridx ),
       .io_bht_update_bits_prediction_bits_target( io_cpu_bht_update_bits_prediction_bits_target ),
       .io_bht_update_bits_prediction_bits_entry( io_cpu_bht_update_bits_prediction_bits_entry ),
       .io_bht_update_bits_prediction_bits_bht_history( io_cpu_bht_update_bits_prediction_bits_bht_history ),
       .io_bht_update_bits_prediction_bits_bht_value( io_cpu_bht_update_bits_prediction_bits_bht_value ),
       .io_bht_update_bits_pc( io_cpu_bht_update_bits_pc ),
       .io_bht_update_bits_taken( io_cpu_bht_update_bits_taken ),
       .io_bht_update_bits_mispredict( io_cpu_bht_update_bits_mispredict ),
       .io_ras_update_valid( io_cpu_ras_update_valid ),
       .io_ras_update_bits_isCall( io_cpu_ras_update_bits_isCall ),
       .io_ras_update_bits_isReturn( io_cpu_ras_update_bits_isReturn ),
       .io_ras_update_bits_returnAddr( io_cpu_ras_update_bits_returnAddr ),
       .io_ras_update_bits_prediction_valid( io_cpu_ras_update_bits_prediction_valid ),
       .io_ras_update_bits_prediction_bits_taken( io_cpu_ras_update_bits_prediction_bits_taken ),
       .io_ras_update_bits_prediction_bits_mask( io_cpu_ras_update_bits_prediction_bits_mask ),
       .io_ras_update_bits_prediction_bits_bridx( io_cpu_ras_update_bits_prediction_bits_bridx ),
       .io_ras_update_bits_prediction_bits_target( io_cpu_ras_update_bits_prediction_bits_target ),
       .io_ras_update_bits_prediction_bits_entry( io_cpu_ras_update_bits_prediction_bits_entry ),
       .io_ras_update_bits_prediction_bits_bht_history( io_cpu_ras_update_bits_prediction_bits_bht_history ),
       .io_ras_update_bits_prediction_bits_bht_value( io_cpu_ras_update_bits_prediction_bits_bht_value ),
       .io_invalidate( T46 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T43 ),
       .io_req_bits_idx( T70 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T39 ),
       .io_resp_ready( Queue_io_enq_ready ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .init( init )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T36 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T35 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_req_bits_store( 1'h0 ),
       .io_resp_miss( tlb_io_resp_miss ),
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( tlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( tlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( tlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( tlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  Queue_9 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( icache_io_resp_valid ),
       //.io_enq_bits_data(  )
       .io_enq_bits_datablock( icache_io_resp_bits_datablock ),
       .io_deq_ready( T0 ),
       .io_deq_valid( Queue_io_deq_valid ),
       //.io_deq_bits_data(  )
       .io_deq_bits_datablock( Queue_io_deq_bits_datablock )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Queue.io_enq_bits_data = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T32) begin
      s1_same_block <= T4;
    end
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T32) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 40'h200;
    end else if(T20) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T32) begin
      s2_valid <= T25;
    end
    if(T52) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T52) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T52) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T52) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T52) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if(T52) begin
      s2_btb_resp_bits_mask <= btb_io_resp_bits_mask;
    end
    if(T52) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T20) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T20) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [1:0] io_req_bits_addr_beat,
    input [25:0] io_req_bits_addr_block,
    input [5:0] io_req_bits_client_xact_id,
    input  io_req_bits_voluntary,
    input [2:0] io_req_bits_r_type,
    input [127:0] io_req_bits_data,
    input [3:0] io_req_bits_way_en,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    //output[3:0] io_meta_read_bits_way_en
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output[3:0] io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[1:0] io_release_bits_addr_beat,
    output[25:0] io_release_bits_addr_block,
    output[5:0] io_release_bits_client_xact_id,
    output io_release_bits_voluntary,
    output[2:0] io_release_bits_r_type,
    output[127:0] io_release_bits_data
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg  req_voluntary;
  wire T2;
  reg [5:0] req_client_xact_id;
  wire[5:0] T3;
  reg [25:0] req_addr_block;
  wire[25:0] T4;
  reg [1:0] beat_cnt;
  wire[1:0] T40;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  reg  r2_data_req_fired;
  wire T41;
  wire T9;
  wire T10;
  reg  r1_data_req_fired;
  wire T42;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg  active;
  wire T43;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [2:0] data_req_cnt;
  wire[2:0] T44;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T45;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[11:0] T33;
  wire[7:0] T34;
  wire[1:0] T35;
  wire[5:0] req_idx;
  reg [3:0] req_way_en;
  wire[3:0] T36;
  wire fire;
  wire T37;
  wire[19:0] T38;
  wire T39;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    req_voluntary = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr_block = {1{$random}};
    beat_cnt = {1{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    data_req_cnt = {1{$random}};
    req_way_en = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_meta_read_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  assign io_release_bits_data = io_data_resp;
  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_voluntary = req_voluntary;
  assign T2 = T1 ? io_req_bits_voluntary : req_voluntary;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T3 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr_block = req_addr_block;
  assign T4 = T1 ? io_req_bits_addr_block : req_addr_block;
  assign io_release_bits_addr_beat = beat_cnt;
  assign T40 = reset ? 2'h0 : T5;
  assign T5 = T7 ? T6 : beat_cnt;
  assign T6 = beat_cnt + 2'h1;
  assign T7 = io_release_ready & io_release_valid;
  assign io_release_valid = T8;
  assign T8 = active & r2_data_req_fired;
  assign T41 = reset ? 1'h0 : T9;
  assign T9 = T18 ? 1'h0 : T10;
  assign T10 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T42 = reset ? 1'h0 : T11;
  assign T11 = T18 ? 1'h0 : T12;
  assign T12 = T14 ? 1'h1 : T13;
  assign T13 = active ? 1'h0 : r1_data_req_fired;
  assign T14 = active & T15;
  assign T15 = T17 & T16;
  assign T16 = io_meta_read_ready & io_meta_read_valid;
  assign T17 = io_data_req_ready & io_data_req_valid;
  assign T18 = T8 & T19;
  assign T19 = io_release_ready ^ 1'h1;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = T1 ? 1'h1 : T21;
  assign T21 = T31 ? T22 : active;
  assign T22 = T24 | T23;
  assign T23 = io_release_ready ^ 1'h1;
  assign T24 = data_req_cnt < 3'h4;
  assign T44 = reset ? 3'h0 : T25;
  assign T25 = T1 ? 3'h0 : T26;
  assign T26 = T18 ? T29 : T27;
  assign T27 = T14 ? T28 : data_req_cnt;
  assign T28 = data_req_cnt + 3'h1;
  assign T29 = data_req_cnt - T45;
  assign T45 = {1'h0, T30};
  assign T30 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign T31 = T8 & T32;
  assign T32 = r1_data_req_fired ^ 1'h1;
  assign io_data_req_bits_addr = T33;
  assign T33 = T34 << 3'h4;
  assign T34 = {req_idx, T35};
  assign T35 = data_req_cnt[1'h1:1'h0];
  assign req_idx = req_addr_block[3'h5:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T36 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T37;
  assign T37 = data_req_cnt < 3'h4;
  assign io_meta_read_bits_tag = T38;
  assign T38 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T39;
  assign T39 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T1) begin
      req_voluntary <= io_req_bits_voluntary;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_addr_block <= io_req_bits_addr_block;
    end
    if(reset) begin
      beat_cnt <= 2'h0;
    end else if(T7) begin
      beat_cnt <= T6;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(T18) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T18) begin
      r1_data_req_fired <= 1'h0;
    end else if(T14) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T31) begin
      active <= T22;
    end
    if(reset) begin
      data_req_cnt <= 3'h0;
    end else if(T1) begin
      data_req_cnt <= 3'h0;
    end else if(T18) begin
      data_req_cnt <= T29;
    end else if(T14) begin
      data_req_cnt <= T28;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_p_type,
    //input [5:0] io_req_bits_client_xact_id
    input  io_rep_ready,
    output io_rep_valid,
    output[1:0] io_rep_bits_addr_beat,
    output[25:0] io_rep_bits_addr_block,
    output[5:0] io_rep_bits_client_xact_id,
    output io_rep_bits_voluntary,
    output[2:0] io_rep_bits_r_type,
    output[127:0] io_rep_bits_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    //output[3:0] io_meta_read_bits_way_en
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[5:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    input [3:0] io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_block_state_state
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg [3:0] way_en;
  wire[3:0] T10;
  wire T11;
  reg [3:0] state;
  wire[3:0] T68;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  wire T29;
  reg [1:0] old_coh_state;
  wire[1:0] T30;
  wire tag_matches;
  wire T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[127:0] reply_data;
  wire[2:0] reply_r_type;
  wire[2:0] T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] miss_coh_state;
  wire T45;
  reg [1:0] req_p_type;
  wire[1:0] T46;
  wire[2:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire T51;
  wire T52;
  wire reply_voluntary;
  wire[5:0] reply_client_xact_id;
  wire[25:0] reply_addr_block;
  reg [25:0] req_addr_block;
  wire[25:0] T53;
  wire[1:0] reply_addr_beat;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[19:0] T62;
  wire[5:0] T69;
  wire T63;
  wire[19:0] T64;
  wire[5:0] T70;
  wire T65;
  wire T66;
  wire T67;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    way_en = {1{$random}};
    state = {1{$random}};
    old_coh_state = {1{$random}};
    req_p_type = {1{$random}};
    req_addr_block = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_meta_read_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T9 | T3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = T6 | T5;
  assign T5 = 3'h2 == io_rep_bits_r_type;
  assign T6 = T8 | T7;
  assign T7 = 3'h1 == io_rep_bits_r_type;
  assign T8 = 3'h0 == io_rep_bits_r_type;
  assign T9 = io_rep_valid ^ 1'h1;
  assign io_wb_req_bits_way_en = way_en;
  assign T10 = T11 ? io_way_en : way_en;
  assign T11 = state == 4'h3;
  assign T68 = reset ? 4'h0 : T12;
  assign T12 = T38 ? 4'h0 : T13;
  assign T13 = T36 ? 4'h8 : T14;
  assign T14 = T35 ? 4'h7 : T15;
  assign T15 = T33 ? T32 : T16;
  assign T16 = T31 ? T27 : T17;
  assign T17 = T25 ? 4'h1 : T18;
  assign T18 = T11 ? 4'h4 : T19;
  assign T19 = T24 ? 4'h3 : T20;
  assign T20 = T23 ? 4'h2 : T21;
  assign T21 = T22 ? 4'h1 : state;
  assign T22 = io_req_ready & io_req_valid;
  assign T23 = io_meta_read_ready & io_meta_read_valid;
  assign T24 = state == 4'h2;
  assign T25 = T11 & T26;
  assign T26 = io_mshr_rdy ^ 1'h1;
  assign T27 = T28 ? 4'h6 : 4'h5;
  assign T28 = tag_matches & T29;
  assign T29 = 2'h3 == old_coh_state;
  assign T30 = T11 ? io_block_state_state : old_coh_state;
  assign tag_matches = way_en != 4'h0;
  assign T31 = state == 4'h4;
  assign T32 = tag_matches ? 4'h8 : 4'h0;
  assign T33 = T34 & io_rep_ready;
  assign T34 = state == 4'h5;
  assign T35 = io_wb_req_ready & io_wb_req_valid;
  assign T36 = T37 & io_wb_req_ready;
  assign T37 = state == 4'h7;
  assign T38 = io_meta_write_ready & io_meta_write_valid;
  assign io_wb_req_bits_data = reply_data;
  assign reply_data = 128'h0;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign reply_r_type = T39;
  assign T39 = T52 ? T50 : T40;
  assign T40 = T49 ? T47 : T41;
  assign T41 = T45 ? T42 : 3'h3;
  assign T42 = T43 ? 3'h2 : 3'h5;
  assign T43 = 2'h3 == T44;
  assign T44 = tag_matches ? old_coh_state : miss_coh_state;
  assign miss_coh_state = 2'h0;
  assign T45 = req_p_type == 2'h2;
  assign T46 = T22 ? io_req_bits_p_type : req_p_type;
  assign T47 = T48 ? 3'h1 : 3'h4;
  assign T48 = 2'h3 == T44;
  assign T49 = req_p_type == 2'h1;
  assign T50 = T51 ? 3'h0 : 3'h3;
  assign T51 = 2'h3 == T44;
  assign T52 = req_p_type == 2'h0;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign reply_voluntary = 1'h0;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign reply_client_xact_id = 6'h0;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign reply_addr_block = req_addr_block;
  assign T53 = T22 ? io_req_bits_addr_block : req_addr_block;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign reply_addr_beat = 2'h0;
  assign io_wb_req_valid = T54;
  assign T54 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T55;
  assign T55 = T56;
  assign T56 = T61 ? 2'h0 : T57;
  assign T57 = T60 ? 2'h1 : T58;
  assign T58 = T59 ? old_coh_state : old_coh_state;
  assign T59 = req_p_type == 2'h2;
  assign T60 = req_p_type == 2'h1;
  assign T61 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T62;
  assign T62 = req_addr_block >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T69;
  assign T69 = req_addr_block[3'h5:1'h0];
  assign io_meta_write_valid = T63;
  assign T63 = state == 4'h8;
  assign io_meta_read_bits_tag = T64;
  assign T64 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = T70;
  assign T70 = req_addr_block[3'h5:1'h0];
  assign io_meta_read_valid = T65;
  assign T65 = state == 4'h1;
  assign io_rep_bits_data = reply_data;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_valid = T66;
  assign T66 = state == 4'h5;
  assign io_req_ready = T67;
  assign T67 = state == 4'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "ProbeUnit should not send releases with data");
    $finish;
  end
// synthesis translate_on
`endif
    if(T11) begin
      way_en <= io_way_en;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T38) begin
      state <= 4'h0;
    end else if(T36) begin
      state <= 4'h8;
    end else if(T35) begin
      state <= 4'h7;
    end else if(T33) begin
      state <= T32;
    end else if(T31) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T11) begin
      state <= 4'h4;
    end else if(T24) begin
      state <= 4'h3;
    end else if(T23) begin
      state <= 4'h2;
    end else if(T22) begin
      state <= 4'h1;
    end
    if(T11) begin
      old_coh_state <= io_block_state_state;
    end
    if(T22) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(T22) begin
      req_addr_block <= io_req_bits_addr_block;
    end
  end
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[19:0] T0;
  wire T1;
  wire[3:0] T2;
  wire[5:0] T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T0;
  assign T0 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T1 = chosen;
  assign io_out_bits_way_en = T2;
  assign T2 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T3;
  assign T3 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T4;
  assign T4 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[1:0] T0;
  wire T1;
  wire[19:0] T2;
  wire[3:0] T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T0;
  assign T0 = T1 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T1 = chosen;
  assign io_out_bits_data_tag = T2;
  assign T2 = T1 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module LockingArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [5:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [127:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [5:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [5:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[5:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  reg [1:0] lockIdx;
  wire[1:0] T67;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T68;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T69;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire[127:0] T22;
  wire[127:0] T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire T29;
  wire T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire T45;
  wire T46;
  wire[25:0] T47;
  wire[25:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid ? 2'h0 : T1;
  assign T1 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T67 = reset ? 2'h2 : T2;
  assign T2 = T7 ? T3 : lockIdx;
  assign T3 = T6 ? 2'h0 : T4;
  assign T4 = T5 ? 2'h1 : 2'h2;
  assign T5 = io_in_1_ready & io_in_1_valid;
  assign T6 = io_in_0_ready & io_in_0_valid;
  assign T7 = T9 & T8;
  assign T8 = locked ^ 1'h1;
  assign T9 = T12 & T10;
  assign T10 = io_out_bits_is_builtin_type & T11;
  assign T11 = 3'h3 == io_out_bits_a_type;
  assign T12 = io_out_valid & io_out_ready;
  assign T68 = reset ? 1'h0 : T13;
  assign T13 = T20 ? 1'h0 : T14;
  assign T14 = T9 ? T15 : locked;
  assign T15 = T16 ^ 1'h1;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T69 = reset ? 2'h0 : T19;
  assign T19 = T9 ? T17 : R18;
  assign T20 = T12 & T21;
  assign T21 = T10 ^ 1'h1;
  assign io_out_bits_data = T22;
  assign T22 = T26 ? io_in_2_bits_data : T23;
  assign T23 = T24 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T24 = T25[1'h0];
  assign T25 = chosen;
  assign T26 = T25[1'h1];
  assign io_out_bits_union = T27;
  assign T27 = T30 ? io_in_2_bits_union : T28;
  assign T28 = T29 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T29 = T25[1'h0];
  assign T30 = T25[1'h1];
  assign io_out_bits_a_type = T31;
  assign T31 = T34 ? io_in_2_bits_a_type : T32;
  assign T32 = T33 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T33 = T25[1'h0];
  assign T34 = T25[1'h1];
  assign io_out_bits_is_builtin_type = T35;
  assign T35 = T38 ? io_in_2_bits_is_builtin_type : T36;
  assign T36 = T37 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T37 = T25[1'h0];
  assign T38 = T25[1'h1];
  assign io_out_bits_addr_beat = T39;
  assign T39 = T42 ? io_in_2_bits_addr_beat : T40;
  assign T40 = T41 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T41 = T25[1'h0];
  assign T42 = T25[1'h1];
  assign io_out_bits_client_xact_id = T43;
  assign T43 = T46 ? io_in_2_bits_client_xact_id : T44;
  assign T44 = T45 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T45 = T25[1'h0];
  assign T46 = T25[1'h1];
  assign io_out_bits_addr_block = T47;
  assign T47 = T50 ? io_in_2_bits_addr_block : T48;
  assign T48 = T49 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T49 = T25[1'h0];
  assign T50 = T25[1'h1];
  assign io_out_valid = T51;
  assign T51 = T54 ? io_in_2_valid : T52;
  assign T52 = T53 ? io_in_1_valid : io_in_0_valid;
  assign T53 = T25[1'h0];
  assign T54 = T25[1'h1];
  assign io_in_0_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = locked ? T57 : 1'h1;
  assign T57 = lockIdx == 2'h0;
  assign io_in_1_ready = T58;
  assign T58 = T59 & io_out_ready;
  assign T59 = locked ? T61 : T60;
  assign T60 = io_in_0_valid ^ 1'h1;
  assign T61 = lockIdx == 2'h1;
  assign io_in_2_ready = T62;
  assign T62 = T63 & io_out_ready;
  assign T63 = locked ? T66 : T64;
  assign T64 = T65 ^ 1'h1;
  assign T65 = io_in_0_valid | io_in_1_valid;
  assign T66 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T7) begin
      lockIdx <= T3;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T20) begin
      locked <= 1'h0;
    end else if(T9) begin
      locked <= T15;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T9) begin
      R18 <= T17;
    end
  end
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [5:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_voluntary,
    input [2:0] io_in_1_bits_r_type,
    input [127:0] io_in_1_bits_data,
    input [3:0] io_in_1_bits_way_en,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [5:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_voluntary,
    input [2:0] io_in_0_bits_r_type,
    input [127:0] io_in_0_bits_data,
    input [3:0] io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[5:0] io_out_bits_client_xact_id,
    output io_out_bits_voluntary,
    output[2:0] io_out_bits_r_type,
    output[127:0] io_out_bits_data,
    output[3:0] io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[3:0] T0;
  wire T1;
  wire[127:0] T2;
  wire[2:0] T3;
  wire T4;
  wire[5:0] T5;
  wire[25:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_way_en = T0;
  assign T0 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_r_type = T3;
  assign T3 = T1 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_voluntary = T4;
  assign T4 = T1 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T6;
  assign T6 = T1 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [39:0] io_in_1_bits_addr,
    input [9:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_kill,
    input  io_in_1_bits_phys,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [9:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_kill,
    input  io_in_0_bits_phys,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[9:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output io_out_bits_kill,
    output io_out_bits_phys,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[4:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire[4:0] T5;
  wire[9:0] T6;
  wire[39:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T0;
  assign T0 = T1 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T1 = chosen;
  assign io_out_bits_phys = T2;
  assign T2 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_kill = T3;
  assign T3 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_bits_typ = T4;
  assign T4 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_cmd = T5;
  assign T5 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T6;
  assign T6 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T7;
  assign T7 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits = T0;
  assign T0 = T1 ? io_in_1_bits : io_in_0_bits;
  assign T1 = chosen;
  assign io_out_valid = T2;
  assign T2 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T3;
  assign T3 = T4 & io_out_ready;
  assign T4 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_20(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [9:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[9:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[64:0] T11;
  reg [64:0] ram [15:0];
  wire[64:0] T12;
  wire[64:0] T13;
  wire[64:0] T14;
  wire[9:0] T15;
  wire[5:0] T16;
  wire[3:0] T17;
  wire[54:0] T18;
  wire[14:0] T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[4:0] T23;
  wire[9:0] T24;
  wire[39:0] T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_phys, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T18 = {io_enq_bits_addr, T19};
  assign T19 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T20;
  assign T20 = T11[3'h5];
  assign io_deq_bits_kill = T21;
  assign T21 = T11[3'h6];
  assign io_deq_bits_typ = T22;
  assign T22 = T11[4'h9:3'h7];
  assign io_deq_bits_cmd = T23;
  assign T23 = T11[4'he:4'ha];
  assign io_deq_bits_tag = T24;
  assign T24 = T11[5'h18:4'hf];
  assign io_deq_bits_addr = T25;
  assign T25 = T11[7'h40:5'h19];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [9:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[5:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    //output[3:0] io_meta_read_bits_way_en
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[9:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[5:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  wire[127:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire T139;
  wire[5:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[5:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[9:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_meta_read_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_voluntary = T139;
  assign T139 = 1'h1;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 6'h0;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 6'h0;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_20 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [9:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[5:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    //output[3:0] io_meta_read_bits_way_en
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[9:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[5:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  wire[127:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire T139;
  wire[5:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[5:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[9:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_meta_read_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_voluntary = T139;
  assign T139 = 1'h1;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 6'h1;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 6'h1;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_20 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module Arbiter_10(
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits = io_in_0_bits;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module Arbiter_11(
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [9:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_nack,
    input  io_in_0_bits_replay,
    input  io_in_0_bits_has_data,
    input [63:0] io_in_0_bits_data_word_bypass,
    input [63:0] io_in_0_bits_store_data,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[9:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output[63:0] io_out_bits_data,
    output io_out_bits_nack,
    output io_out_bits_replay,
    output io_out_bits_has_data,
    output[63:0] io_out_bits_data_word_bypass,
    output[63:0] io_out_bits_store_data,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_nack = io_in_0_bits_nack;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module IOMSHR(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [9:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_acquire_ready,
    output io_acquire_valid,
    output[25:0] io_acquire_bits_addr_block,
    output[5:0] io_acquire_bits_client_xact_id,
    output[1:0] io_acquire_bits_addr_beat,
    output io_acquire_bits_is_builtin_type,
    output[2:0] io_acquire_bits_a_type,
    output[16:0] io_acquire_bits_union,
    output[127:0] io_acquire_bits_data,
    input  io_grant_valid,
    input [1:0] io_grant_bits_addr_beat,
    input [5:0] io_grant_bits_client_xact_id,
    input [3:0] io_grant_bits_manager_xact_id,
    input  io_grant_bits_is_builtin_type,
    input [3:0] io_grant_bits_g_type,
    input [127:0] io_grant_bits_data,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[9:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    //output[63:0] io_resp_bits_data_word_bypass
    output[63:0] io_resp_bits_store_data
);

  reg [63:0] req_data;
  wire[63:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg [4:0] req_cmd;
  wire[4:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] T141;
  wire req_cmd_sc;
  wire[63:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire[7:0] T16;
  wire[63:0] T17;
  wire[15:0] T18;
  wire[15:0] T19;
  wire[63:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  reg [63:0] grant_word;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[127:0] T25;
  wire[6:0] T26;
  wire T27;
  reg [39:0] req_addr;
  wire[39:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg [1:0] state;
  wire[1:0] T142;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T143;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  reg [2:0] req_typ;
  wire[2:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[15:0] T62;
  wire T63;
  wire[47:0] T64;
  wire[47:0] T65;
  wire[47:0] T66;
  wire[47:0] T144;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire[55:0] T72;
  wire[55:0] T73;
  wire[55:0] T74;
  wire[55:0] T145;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [9:0] req_tag;
  wire[9:0] T79;
  wire T80;
  wire[127:0] T81;
  wire[127:0] put_acquire_data;
  wire[127:0] beat_data;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[31:0] T86;
  wire T87;
  wire[1:0] T88;
  wire[63:0] T89;
  wire[31:0] T90;
  wire[15:0] T91;
  wire T92;
  wire[63:0] T93;
  wire[31:0] T94;
  wire[15:0] T95;
  wire[7:0] T96;
  wire T97;
  wire[127:0] get_acquire_data;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[16:0] T107;
  wire[16:0] put_acquire_union;
  wire[16:0] T146;
  wire[23:0] T108;
  wire[22:0] beat_mask;
  wire[3:0] T109;
  wire beat_offset;
  wire[7:0] T110;
  wire[3:0] T111;
  wire[3:0] T112;
  wire[1:0] T113;
  wire[1:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire T129;
  wire[3:0] T130;
  wire T131;
  wire[16:0] get_acquire_union;
  wire[16:0] T147;
  wire[12:0] T132;
  wire[6:0] T133;
  wire[3:0] addr_byte;
  wire[2:0] T134;
  wire[2:0] put_acquire_a_type;
  wire[2:0] get_acquire_a_type;
  wire T135;
  wire put_acquire_is_builtin_type;
  wire get_acquire_is_builtin_type;
  wire[1:0] T136;
  wire[1:0] put_acquire_addr_beat;
  wire[1:0] addr_beat;
  wire[1:0] get_acquire_addr_beat;
  wire[5:0] T137;
  wire[5:0] put_acquire_client_xact_id;
  wire[5:0] get_acquire_client_xact_id;
  wire[25:0] T138;
  wire[25:0] put_acquire_addr_block;
  wire[25:0] addr_block;
  wire[25:0] get_acquire_addr_block;
  wire T139;
  wire T140;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_data = {2{$random}};
    req_cmd = {1{$random}};
    grant_word = {2{$random}};
    req_addr = {2{$random}};
    state = {1{$random}};
    req_typ = {1{$random}};
    req_tag = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_resp_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  assign io_resp_bits_store_data = req_data;
  assign T0 = T1 ? io_req_bits_data : req_data;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_has_data = T2;
  assign T2 = T7 | T3;
  assign T3 = T6 | T4;
  assign T4 = req_cmd == 5'h4;
  assign T5 = T1 ? io_req_bits_cmd : req_cmd;
  assign T6 = req_cmd[2'h3];
  assign T7 = T9 | T8;
  assign T8 = req_cmd == 5'h7;
  assign T9 = T11 | T10;
  assign T10 = req_cmd == 5'h6;
  assign T11 = req_cmd == 5'h0;
  assign io_resp_bits_replay = io_resp_valid;
  assign io_resp_bits_nack = 1'h0;
  assign io_resp_bits_data = T12;
  assign T12 = T13 | T141;
  assign T141 = {63'h0, req_cmd_sc};
  assign req_cmd_sc = req_cmd == 5'h7;
  assign T13 = {T72, T14};
  assign T14 = req_cmd_sc ? 8'h0 : T15;
  assign T15 = T71 ? T70 : T16;
  assign T16 = T17[3'h7:1'h0];
  assign T17 = {T64, T18};
  assign T18 = T63 ? T62 : T19;
  assign T19 = T20[4'hf:1'h0];
  assign T20 = {T52, T21};
  assign T21 = T51 ? T50 : T22;
  assign T22 = grant_word[5'h1f:1'h0];
  assign T23 = T29 ? T24 : grant_word;
  assign T24 = T25[6'h3f:1'h0];
  assign T25 = io_grant_bits_data >> T26;
  assign T26 = {T27, 6'h0};
  assign T27 = req_addr[2'h3];
  assign T28 = T1 ? io_req_bits_addr : req_addr;
  assign T29 = T39 & T30;
  assign T30 = T34 | T31;
  assign T31 = T33 | T32;
  assign T32 = req_cmd == 5'h4;
  assign T33 = req_cmd[2'h3];
  assign T34 = T36 | T35;
  assign T35 = req_cmd == 5'h7;
  assign T36 = T38 | T37;
  assign T37 = req_cmd == 5'h6;
  assign T38 = req_cmd == 5'h0;
  assign T39 = T40 & io_grant_valid;
  assign T40 = state == 2'h2;
  assign T142 = reset ? 2'h0 : T41;
  assign T41 = T49 ? 2'h0 : T42;
  assign T42 = T47 ? 2'h0 : T43;
  assign T43 = T29 ? 2'h3 : T44;
  assign T44 = T46 ? 2'h2 : T45;
  assign T45 = T1 ? 2'h1 : state;
  assign T46 = io_acquire_ready & io_acquire_valid;
  assign T47 = T39 & T48;
  assign T48 = T30 ^ 1'h1;
  assign T49 = io_resp_ready & io_resp_valid;
  assign T50 = grant_word[6'h3f:6'h20];
  assign T51 = req_addr[2'h2];
  assign T52 = T60 ? T54 : T53;
  assign T53 = grant_word[6'h3f:6'h20];
  assign T54 = 32'h0 - T143;
  assign T143 = {31'h0, T55};
  assign T55 = T57 & T56;
  assign T56 = T21[5'h1f];
  assign T57 = $signed(1'h0) <= $signed(T58);
  assign T58 = req_typ;
  assign T59 = T1 ? io_req_bits_typ : req_typ;
  assign T60 = T61 == 2'h2;
  assign T61 = req_typ[1'h1:1'h0];
  assign T62 = T20[5'h1f:5'h10];
  assign T63 = req_addr[1'h1];
  assign T64 = T69 ? T66 : T65;
  assign T65 = T20[6'h3f:5'h10];
  assign T66 = 48'h0 - T144;
  assign T144 = {47'h0, T67};
  assign T67 = T57 & T68;
  assign T68 = T18[4'hf];
  assign T69 = T61 == 2'h1;
  assign T70 = T17[4'hf:4'h8];
  assign T71 = req_addr[1'h0];
  assign T72 = T77 ? T74 : T73;
  assign T73 = T17[6'h3f:4'h8];
  assign T74 = 56'h0 - T145;
  assign T145 = {55'h0, T75};
  assign T75 = T57 & T76;
  assign T76 = T14[3'h7];
  assign T77 = T78 | req_cmd_sc;
  assign T78 = T61 == 2'h0;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_tag = req_tag;
  assign T79 = T1 ? io_req_bits_tag : req_tag;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_valid = T80;
  assign T80 = state == 2'h3;
  assign io_acquire_bits_data = T81;
  assign T81 = T98 ? get_acquire_data : put_acquire_data;
  assign put_acquire_data = beat_data;
  assign beat_data = {T82, T82};
  assign T82 = T97 ? T93 : T83;
  assign T83 = T92 ? T89 : T84;
  assign T84 = T87 ? T85 : req_data;
  assign T85 = {T86, T86};
  assign T86 = req_data[5'h1f:1'h0];
  assign T87 = T88 == 2'h2;
  assign T88 = req_typ[1'h1:1'h0];
  assign T89 = {T90, T90};
  assign T90 = {T91, T91};
  assign T91 = req_data[4'hf:1'h0];
  assign T92 = T88 == 2'h1;
  assign T93 = {T94, T94};
  assign T94 = {T95, T95};
  assign T95 = {T96, T96};
  assign T96 = req_data[3'h7:1'h0];
  assign T97 = T88 == 2'h0;
  assign get_acquire_data = 128'h0;
  assign T98 = T102 | T99;
  assign T99 = T101 | T100;
  assign T100 = req_cmd == 5'h4;
  assign T101 = req_cmd[2'h3];
  assign T102 = T104 | T103;
  assign T103 = req_cmd == 5'h7;
  assign T104 = T106 | T105;
  assign T105 = req_cmd == 5'h6;
  assign T106 = req_cmd == 5'h0;
  assign io_acquire_bits_union = T107;
  assign T107 = T98 ? get_acquire_union : put_acquire_union;
  assign put_acquire_union = T146;
  assign T146 = T108[5'h10:1'h0];
  assign T108 = {beat_mask, 1'h0};
  assign beat_mask = T110 << T109;
  assign T109 = {beat_offset, 3'h0};
  assign beat_offset = req_addr[2'h3];
  assign T110 = {T127, T111};
  assign T111 = T126 ? 4'h0 : T112;
  assign T112 = {T121, T113};
  assign T113 = T120 ? 2'h0 : T114;
  assign T114 = {T117, T115};
  assign T115 = T116 == 1'h0;
  assign T116 = req_addr[1'h0];
  assign T117 = T119 | T118;
  assign T118 = 2'h1 <= T88;
  assign T119 = req_addr[1'h0];
  assign T120 = req_addr[1'h1];
  assign T121 = T124 | T122;
  assign T122 = T123 ? 2'h3 : 2'h0;
  assign T123 = 2'h2 <= T88;
  assign T124 = T125 ? T114 : 2'h0;
  assign T125 = req_addr[1'h1];
  assign T126 = req_addr[2'h2];
  assign T127 = T130 | T128;
  assign T128 = T129 ? 4'hf : 4'h0;
  assign T129 = 2'h3 <= T88;
  assign T130 = T131 ? T112 : 4'h0;
  assign T131 = req_addr[2'h2];
  assign get_acquire_union = T147;
  assign T147 = {4'h0, T132};
  assign T132 = {T133, 6'h0};
  assign T133 = {addr_byte, req_typ};
  assign addr_byte = req_addr[2'h3:1'h0];
  assign io_acquire_bits_a_type = T134;
  assign T134 = T98 ? get_acquire_a_type : put_acquire_a_type;
  assign put_acquire_a_type = 3'h2;
  assign get_acquire_a_type = 3'h0;
  assign io_acquire_bits_is_builtin_type = T135;
  assign T135 = T98 ? get_acquire_is_builtin_type : put_acquire_is_builtin_type;
  assign put_acquire_is_builtin_type = 1'h1;
  assign get_acquire_is_builtin_type = 1'h1;
  assign io_acquire_bits_addr_beat = T136;
  assign T136 = T98 ? get_acquire_addr_beat : put_acquire_addr_beat;
  assign put_acquire_addr_beat = addr_beat;
  assign addr_beat = req_addr[3'h5:3'h4];
  assign get_acquire_addr_beat = addr_beat;
  assign io_acquire_bits_client_xact_id = T137;
  assign T137 = T98 ? get_acquire_client_xact_id : put_acquire_client_xact_id;
  assign put_acquire_client_xact_id = 6'h2;
  assign get_acquire_client_xact_id = 6'h2;
  assign io_acquire_bits_addr_block = T138;
  assign T138 = T98 ? get_acquire_addr_block : put_acquire_addr_block;
  assign put_acquire_addr_block = addr_block;
  assign addr_block = req_addr[5'h1f:3'h6];
  assign get_acquire_addr_block = addr_block;
  assign io_acquire_valid = T139;
  assign T139 = state == 2'h1;
  assign io_req_ready = T140;
  assign T140 = state == 2'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_data <= io_req_bits_data;
    end
    if(T1) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T29) begin
      grant_word <= T24;
    end
    if(T1) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T49) begin
      state <= 2'h0;
    end else if(T47) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= 2'h3;
    end else if(T46) begin
      state <= 2'h2;
    end else if(T1) begin
      state <= 2'h1;
    end
    if(T1) begin
      req_typ <= io_req_bits_typ;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [9:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[9:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    output[63:0] io_resp_bits_data_word_bypass,
    output[63:0] io_resp_bits_store_data,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[5:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output[3:0] io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[3:0] io_meta_read_bits_way_en,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[9:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[5:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output[3:0] io_wb_req_bits_way_en,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire cacheable;
  wire T4;
  wire T5;
  wire[4:0] T111;
  wire[4:0] T112;
  wire[4:0] T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire[4:0] T116;
  wire[4:0] T117;
  wire[4:0] T118;
  wire[4:0] T119;
  wire[4:0] T120;
  wire[4:0] T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire[4:0] T124;
  wire[4:0] T125;
  wire[4:0] T126;
  wire T127;
  wire[16:0] T6;
  wire[16:0] T7;
  reg [16:0] sdq_val;
  wire[16:0] T128;
  wire[31:0] T129;
  wire[31:0] T8;
  wire[31:0] T130;
  wire[31:0] T9;
  wire[31:0] T131;
  wire[16:0] T10;
  wire[16:0] T11;
  wire[16:0] T132;
  wire sdq_enq;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[16:0] T23;
  wire[16:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[31:0] T57;
  wire[31:0] T58;
  wire[31:0] T59;
  wire[31:0] T133;
  wire[16:0] T60;
  wire[16:0] T134;
  wire free_sdq;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire[31:0] T69;
  wire[31:0] T135;
  wire T70;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T71;
  wire tag_match;
  wire[27:0] T72;
  wire[27:0] T151;
  wire[19:0] T73;
  wire[19:0] T74;
  wire[19:0] tagList_1;
  wire idxMatch_1;
  wire[19:0] T75;
  wire[19:0] tagList_0;
  wire idxMatch_0;
  wire T76;
  wire sdq_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire idx_match;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[63:0] T96;
  reg [63:0] sdq [16:0];
  wire[63:0] T97;
  wire T98;
  wire T99;
  wire[4:0] T100;
  reg [4:0] R101;
  wire[4:0] T102;
  wire[11:0] T103;
  wire[11:0] refillMux_0_addr;
  wire[11:0] refillMux_1_addr;
  wire T104;
  wire T152;
  wire[3:0] T105;
  wire[3:0] refillMux_0_way_en;
  wire[3:0] refillMux_1_way_en;
  wire T106;
  wire T107;
  wire T108;
  wire pri_rdy;
  wire T109;
  wire sec_rdy;
  wire T110;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire[3:0] meta_read_arb_io_out_bits_way_en;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire[3:0] meta_write_arb_io_out_bits_way_en;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_2_ready;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr_block;
  wire[5:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[1:0] mem_req_arb_io_out_bits_addr_beat;
  wire mem_req_arb_io_out_bits_is_builtin_type;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[16:0] mem_req_arb_io_out_bits_union;
  wire[127:0] mem_req_arb_io_out_bits_data;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[1:0] wb_req_arb_io_out_bits_addr_beat;
  wire[25:0] wb_req_arb_io_out_bits_addr_block;
  wire[5:0] wb_req_arb_io_out_bits_client_xact_id;
  wire wb_req_arb_io_out_bits_voluntary;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire[127:0] wb_req_arb_io_out_bits_data;
  wire[3:0] wb_req_arb_io_out_bits_way_en;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire[39:0] replay_arb_io_out_bits_addr;
  wire[9:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_bits_phys;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire mmio_alloc_arb_io_in_0_ready;
  wire resp_arb_io_in_0_ready;
  wire resp_arb_io_out_valid;
  wire[39:0] resp_arb_io_out_bits_addr;
  wire[9:0] resp_arb_io_out_bits_tag;
  wire[4:0] resp_arb_io_out_bits_cmd;
  wire[2:0] resp_arb_io_out_bits_typ;
  wire[63:0] resp_arb_io_out_bits_data;
  wire resp_arb_io_out_bits_nack;
  wire resp_arb_io_out_bits_replay;
  wire resp_arb_io_out_bits_has_data;
  wire[63:0] resp_arb_io_out_bits_data_word_bypass;
  wire[63:0] resp_arb_io_out_bits_store_data;
  wire IOMSHR_io_req_ready;
  wire IOMSHR_io_acquire_valid;
  wire[25:0] IOMSHR_io_acquire_bits_addr_block;
  wire[5:0] IOMSHR_io_acquire_bits_client_xact_id;
  wire[1:0] IOMSHR_io_acquire_bits_addr_beat;
  wire IOMSHR_io_acquire_bits_is_builtin_type;
  wire[2:0] IOMSHR_io_acquire_bits_a_type;
  wire[16:0] IOMSHR_io_acquire_bits_union;
  wire[127:0] IOMSHR_io_acquire_bits_data;
  wire IOMSHR_io_resp_valid;
  wire[39:0] IOMSHR_io_resp_bits_addr;
  wire[9:0] IOMSHR_io_resp_bits_tag;
  wire[4:0] IOMSHR_io_resp_bits_cmd;
  wire[2:0] IOMSHR_io_resp_bits_typ;
  wire[63:0] IOMSHR_io_resp_bits_data;
  wire IOMSHR_io_resp_bits_nack;
  wire IOMSHR_io_resp_bits_replay;
  wire IOMSHR_io_resp_bits_has_data;
  wire[63:0] IOMSHR_io_resp_bits_store_data;
  wire MSHR_io_req_pri_rdy;
  wire MSHR_io_req_sec_rdy;
  wire MSHR_io_idx_match;
  wire[19:0] MSHR_io_tag;
  wire MSHR_io_mem_req_valid;
  wire[25:0] MSHR_io_mem_req_bits_addr_block;
  wire[5:0] MSHR_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_io_mem_req_bits_addr_beat;
  wire MSHR_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_io_mem_req_bits_a_type;
  wire[16:0] MSHR_io_mem_req_bits_union;
  wire[127:0] MSHR_io_mem_req_bits_data;
  wire[3:0] MSHR_io_refill_way_en;
  wire[11:0] MSHR_io_refill_addr;
  wire MSHR_io_meta_read_valid;
  wire[5:0] MSHR_io_meta_read_bits_idx;
  wire[19:0] MSHR_io_meta_read_bits_tag;
  wire MSHR_io_meta_write_valid;
  wire[5:0] MSHR_io_meta_write_bits_idx;
  wire[3:0] MSHR_io_meta_write_bits_way_en;
  wire[19:0] MSHR_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_io_meta_write_bits_data_coh_state;
  wire MSHR_io_replay_valid;
  wire[39:0] MSHR_io_replay_bits_addr;
  wire[9:0] MSHR_io_replay_bits_tag;
  wire[4:0] MSHR_io_replay_bits_cmd;
  wire[2:0] MSHR_io_replay_bits_typ;
  wire MSHR_io_replay_bits_kill;
  wire MSHR_io_replay_bits_phys;
  wire[4:0] MSHR_io_replay_bits_sdq_id;
  wire MSHR_io_wb_req_valid;
  wire[1:0] MSHR_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_io_wb_req_bits_addr_block;
  wire[5:0] MSHR_io_wb_req_bits_client_xact_id;
  wire MSHR_io_wb_req_bits_voluntary;
  wire[2:0] MSHR_io_wb_req_bits_r_type;
  wire[127:0] MSHR_io_wb_req_bits_data;
  wire[3:0] MSHR_io_wb_req_bits_way_en;
  wire MSHR_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[19:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr_block;
  wire[5:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_1_io_mem_req_bits_addr_beat;
  wire MSHR_1_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[16:0] MSHR_1_io_mem_req_bits_union;
  wire[127:0] MSHR_1_io_mem_req_bits_data;
  wire[3:0] MSHR_1_io_refill_way_en;
  wire[11:0] MSHR_1_io_refill_addr;
  wire MSHR_1_io_meta_read_valid;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire[3:0] MSHR_1_io_meta_write_bits_way_en;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire[39:0] MSHR_1_io_replay_bits_addr;
  wire[9:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_bits_phys;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_wb_req_valid;
  wire[1:0] MSHR_1_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_1_io_wb_req_bits_addr_block;
  wire[5:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire MSHR_1_io_wb_req_bits_voluntary;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire[127:0] MSHR_1_io_wb_req_bits_data;
  wire[3:0] MSHR_1_io_wb_req_bits_way_en;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R101 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_grant_valid & T1;
  assign T1 = io_mem_grant_bits_client_xact_id == 6'h2;
  assign T2 = io_req_valid & T3;
  assign T3 = cacheable ^ 1'h1;
  assign cacheable = io_req_bits_addr < 40'h40000000;
  assign T4 = io_mem_grant_valid & T5;
  assign T5 = io_mem_grant_bits_client_xact_id == 6'h1;
  assign T111 = T150 ? 1'h0 : T112;
  assign T112 = T149 ? 1'h1 : T113;
  assign T113 = T148 ? 2'h2 : T114;
  assign T114 = T147 ? 2'h3 : T115;
  assign T115 = T146 ? 3'h4 : T116;
  assign T116 = T145 ? 3'h5 : T117;
  assign T117 = T144 ? 3'h6 : T118;
  assign T118 = T143 ? 3'h7 : T119;
  assign T119 = T142 ? 4'h8 : T120;
  assign T120 = T141 ? 4'h9 : T121;
  assign T121 = T140 ? 4'ha : T122;
  assign T122 = T139 ? 4'hb : T123;
  assign T123 = T138 ? 4'hc : T124;
  assign T124 = T137 ? 4'hd : T125;
  assign T125 = T136 ? 4'he : T126;
  assign T126 = T127 ? 4'hf : 5'h10;
  assign T127 = T6[4'hf];
  assign T6 = ~ T7;
  assign T7 = sdq_val;
  assign T128 = T129[5'h10:1'h0];
  assign T129 = reset ? 32'h0 : T8;
  assign T8 = T70 ? T9 : T130;
  assign T130 = {15'h0, sdq_val};
  assign T9 = T57 | T131;
  assign T131 = {15'h0, T10};
  assign T10 = T21 & T11;
  assign T11 = 17'h0 - T132;
  assign T132 = {16'h0, sdq_enq};
  assign sdq_enq = T19 & T12;
  assign T12 = T16 | T13;
  assign T13 = T15 | T14;
  assign T14 = io_req_bits_cmd == 5'h4;
  assign T15 = io_req_bits_cmd[2'h3];
  assign T16 = T18 | T17;
  assign T17 = io_req_bits_cmd == 5'h7;
  assign T18 = io_req_bits_cmd == 5'h1;
  assign T19 = T20 & cacheable;
  assign T20 = io_req_valid & io_req_ready;
  assign T21 = T56 ? 17'h1 : T22;
  assign T22 = T55 ? 17'h2 : T23;
  assign T23 = T54 ? 17'h4 : T24;
  assign T24 = T53 ? 17'h8 : T25;
  assign T25 = T52 ? 17'h10 : T26;
  assign T26 = T51 ? 17'h20 : T27;
  assign T27 = T50 ? 17'h40 : T28;
  assign T28 = T49 ? 17'h80 : T29;
  assign T29 = T48 ? 17'h100 : T30;
  assign T30 = T47 ? 17'h200 : T31;
  assign T31 = T46 ? 17'h400 : T32;
  assign T32 = T45 ? 17'h800 : T33;
  assign T33 = T44 ? 17'h1000 : T34;
  assign T34 = T43 ? 17'h2000 : T35;
  assign T35 = T42 ? 17'h4000 : T36;
  assign T36 = T41 ? 17'h8000 : T37;
  assign T37 = T38 ? 17'h10000 : 17'h0;
  assign T38 = T39[5'h10];
  assign T39 = ~ T40;
  assign T40 = sdq_val;
  assign T41 = T39[4'hf];
  assign T42 = T39[4'he];
  assign T43 = T39[4'hd];
  assign T44 = T39[4'hc];
  assign T45 = T39[4'hb];
  assign T46 = T39[4'ha];
  assign T47 = T39[4'h9];
  assign T48 = T39[4'h8];
  assign T49 = T39[3'h7];
  assign T50 = T39[3'h6];
  assign T51 = T39[3'h5];
  assign T52 = T39[3'h4];
  assign T53 = T39[2'h3];
  assign T54 = T39[2'h2];
  assign T55 = T39[1'h1];
  assign T56 = T39[1'h0];
  assign T57 = T135 & T58;
  assign T58 = ~ T59;
  assign T59 = T69 & T133;
  assign T133 = {15'h0, T60};
  assign T60 = 17'h0 - T134;
  assign T134 = {16'h0, free_sdq};
  assign free_sdq = T68 & T61;
  assign T61 = T65 | T62;
  assign T62 = T64 | T63;
  assign T63 = io_replay_bits_cmd == 5'h4;
  assign T64 = io_replay_bits_cmd[2'h3];
  assign T65 = T67 | T66;
  assign T66 = io_replay_bits_cmd == 5'h7;
  assign T67 = io_replay_bits_cmd == 5'h1;
  assign T68 = io_replay_ready & io_replay_valid;
  assign T69 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T135 = {15'h0, sdq_val};
  assign T70 = io_replay_valid | sdq_enq;
  assign T136 = T6[4'he];
  assign T137 = T6[4'hd];
  assign T138 = T6[4'hc];
  assign T139 = T6[4'hb];
  assign T140 = T6[4'ha];
  assign T141 = T6[4'h9];
  assign T142 = T6[4'h8];
  assign T143 = T6[3'h7];
  assign T144 = T6[3'h6];
  assign T145 = T6[3'h5];
  assign T146 = T6[3'h4];
  assign T147 = T6[2'h3];
  assign T148 = T6[2'h2];
  assign T149 = T6[1'h1];
  assign T150 = T6[1'h0];
  assign T71 = T76 & tag_match;
  assign tag_match = T151 == T72;
  assign T72 = io_req_bits_addr >> 4'hc;
  assign T151 = {8'h0, T73};
  assign T73 = T75 | T74;
  assign T74 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T75 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_io_tag;
  assign idxMatch_0 = MSHR_io_idx_match;
  assign T76 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T77 ^ 1'h1;
  assign T77 = sdq_val == 17'h1ffff;
  assign T78 = io_mem_grant_valid & T79;
  assign T79 = io_mem_grant_bits_client_xact_id == 6'h0;
  assign T80 = T81 & tag_match;
  assign T81 = io_req_valid & sdq_rdy;
  assign T82 = T84 & T83;
  assign T83 = idx_match ^ 1'h1;
  assign idx_match = MSHR_io_idx_match | MSHR_1_io_idx_match;
  assign T84 = T85 & cacheable;
  assign T85 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T86;
  assign T86 = T91 ? 1'h0 : T87;
  assign T87 = T90 ? 1'h0 : T88;
  assign T88 = T89 == 1'h0;
  assign T89 = MSHR_io_req_pri_rdy ^ 1'h1;
  assign T90 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign T91 = IOMSHR_io_req_ready ^ 1'h1;
  assign io_probe_rdy = T92;
  assign T92 = T95 ? 1'h0 : T93;
  assign T93 = T94 == 1'h0;
  assign T94 = MSHR_io_probe_rdy ^ 1'h1;
  assign T95 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_replay_bits_data = T96;
  assign T96 = sdq[R101];
  assign T98 = sdq_enq & T99;
  assign T99 = T100 < 5'h11;
  assign T100 = T111;
  assign T102 = free_sdq ? replay_arb_io_out_bits_sdq_id : R101;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_way_en = meta_read_arb_io_out_bits_way_en;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_refill_addr = T103;
  assign T103 = T104 ? refillMux_1_addr : refillMux_0_addr;
  assign refillMux_0_addr = MSHR_io_refill_addr;
  assign refillMux_1_addr = MSHR_1_io_refill_addr;
  assign T104 = T152;
  assign T152 = io_mem_grant_bits_client_xact_id[1'h0];
  assign io_refill_way_en = T105;
  assign T105 = T104 ? refillMux_1_way_en : refillMux_0_way_en;
  assign refillMux_0_way_en = MSHR_io_refill_way_en;
  assign refillMux_1_way_en = MSHR_1_io_refill_way_en;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_nack = resp_arb_io_out_bits_nack;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_req_ready = T106;
  assign T106 = T110 ? IOMSHR_io_req_ready : T107;
  assign T107 = T108 & sdq_rdy;
  assign T108 = idx_match ? T109 : pri_rdy;
  assign pri_rdy = MSHR_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T109 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  assign T110 = cacheable ^ 1'h1;
  Arbiter_7 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       //.io_in_1_bits_way_en(  )
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_read_bits_idx ),
       //.io_in_0_bits_way_en(  )
       .io_in_0_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_read_arb_io_out_bits_way_en ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign meta_read_arb.io_in_1_bits_way_en = {1{$random}};
    assign meta_read_arb.io_in_0_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  LockingArbiter_1 mem_req_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( mem_req_arb_io_in_2_ready ),
       .io_in_2_valid( IOMSHR_io_acquire_valid ),
       .io_in_2_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_in_2_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_in_2_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_in_2_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_mem_req_valid ),
       .io_in_0_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_in_0_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_in_0_bits_union( MSHR_io_mem_req_bits_union ),
       .io_in_0_bits_data( MSHR_io_mem_req_bits_data ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr_block( mem_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( mem_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( mem_req_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_union( mem_req_arb_io_out_bits_union ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_1_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_in_0_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_in_0_bits_data( MSHR_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_addr_beat( wb_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wb_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( wb_req_arb_io_out_bits_voluntary ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type ),
       .io_out_bits_data( wb_req_arb_io_out_bits_data ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en )
       //.io_chosen(  )
  );
  Arbiter_8 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_replay_valid ),
       .io_in_0_bits_addr( MSHR_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_in_0_bits_typ( MSHR_io_replay_bits_typ ),
       .io_in_0_bits_kill( MSHR_io_replay_bits_kill ),
       .io_in_0_bits_phys( MSHR_io_replay_bits_phys ),
       .io_in_0_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_9 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T82 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  MSHR_0 MSHR(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_io_req_pri_rdy ),
       .io_req_sec_val( T80 ),
       .io_req_sec_rdy( MSHR_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T111 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_io_idx_match ),
       .io_tag( MSHR_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_io_refill_way_en ),
       .io_refill_addr( MSHR_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_io_meta_read_bits_idx ),
       //.io_meta_read_bits_way_en(  )
       .io_meta_read_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_io_replay_valid ),
       .io_replay_bits_addr( MSHR_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T78 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( MSHR_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_io_probe_rdy )
  );
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T71 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T111 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_1_io_refill_way_en ),
       .io_refill_addr( MSHR_1_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       //.io_meta_read_bits_way_en(  )
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T4 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  Arbiter_10 mmio_alloc_arb(
       .io_in_0_ready( mmio_alloc_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_req_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T2 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign mmio_alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_11 resp_arb(
       .io_in_0_ready( resp_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_resp_valid ),
       .io_in_0_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_in_0_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_in_0_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_in_0_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_in_0_bits_data( IOMSHR_io_resp_bits_data ),
       .io_in_0_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_in_0_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_in_0_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_in_0_bits_data_word_bypass(  )
       .io_in_0_bits_store_data( IOMSHR_io_resp_bits_store_data ),
       .io_out_ready( io_resp_ready ),
       .io_out_valid( resp_arb_io_out_valid ),
       .io_out_bits_addr( resp_arb_io_out_bits_addr ),
       .io_out_bits_tag( resp_arb_io_out_bits_tag ),
       .io_out_bits_cmd( resp_arb_io_out_bits_cmd ),
       .io_out_bits_typ( resp_arb_io_out_bits_typ ),
       .io_out_bits_data( resp_arb_io_out_bits_data ),
       .io_out_bits_nack( resp_arb_io_out_bits_nack ),
       .io_out_bits_replay( resp_arb_io_out_bits_replay ),
       .io_out_bits_has_data( resp_arb_io_out_bits_has_data ),
       .io_out_bits_data_word_bypass( resp_arb_io_out_bits_data_word_bypass ),
       .io_out_bits_store_data( resp_arb_io_out_bits_store_data )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign resp_arb.io_in_0_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  IOMSHR IOMSHR(.clk(clk), .reset(reset),
       .io_req_ready( IOMSHR_io_req_ready ),
       .io_req_valid( mmio_alloc_arb_io_in_0_ready ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_data( io_req_bits_data ),
       .io_acquire_ready( mem_req_arb_io_in_2_ready ),
       .io_acquire_valid( IOMSHR_io_acquire_valid ),
       .io_acquire_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_acquire_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_acquire_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_acquire_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_acquire_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_acquire_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_acquire_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_grant_valid( T0 ),
       .io_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_grant_bits_data( io_mem_grant_bits_data ),
       .io_resp_ready( resp_arb_io_in_0_ready ),
       .io_resp_valid( IOMSHR_io_resp_valid ),
       .io_resp_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_resp_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_resp_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_resp_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_resp_bits_data( IOMSHR_io_resp_bits_data ),
       .io_resp_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_resp_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_resp_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( IOMSHR_io_resp_bits_store_data )
  );

  always @(posedge clk) begin
    sdq_val <= T128;
    if (T98)
      sdq[T111] <= io_req_bits_data;
    if(free_sdq) begin
      R101 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    input [3:0] io_read_bits_way_en,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input [3:0] io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_3_tag,
    output[1:0] io_resp_3_coh_state,
    output[19:0] io_resp_2_tag,
    output[1:0] io_resp_2_coh_state,
    output[19:0] io_resp_1_tag,
    output[1:0] io_resp_1_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state,
    input  init
);

  wire[1:0] T0;
  wire[87:0] T1;
  wire[87:0] T2;
  wire[43:0] T3;
  wire[21:0] T4;
  wire[87:0] T5;
  wire[87:0] T7;
  wire[87:0] T8;
  wire[87:0] T9;
  wire[43:0] T10;
  wire[21:0] T11;
  wire[21:0] T50;
  wire T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T51;
  wire[6:0] T15;
  wire[6:0] T16;
  wire[21:0] T17;
  wire[21:0] T52;
  wire T18;
  wire[43:0] T19;
  wire[21:0] T20;
  wire[21:0] T53;
  wire T21;
  wire[21:0] T22;
  wire[21:0] T54;
  wire T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[43:0] T26;
  wire[21:0] wdata;
  wire[21:0] T27;
  wire[1:0] T28;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T29;
  wire[19:0] T30;
  wire[19:0] rstVal_tag;
  wire[43:0] T31;
  wire T32;
  wire[5:0] T55;
  wire[6:0] waddr;
  wire[6:0] T56;
  reg [5:0] R33;
  wire[5:0] T34;
  wire[21:0] T35;
  wire[43:0] T36;
  wire[21:0] T37;
  wire[21:0] T38;
  wire[19:0] T39;
  wire[1:0] T40;
  wire[19:0] T41;
  wire[1:0] T42;
  wire[19:0] T43;
  wire[1:0] T44;
  wire[19:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R33 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = T2;
  assign T2 = {T36, T3};
  assign T3 = {T35, T4};
  assign T4 = T5[5'h15:1'h0];
  MetadataArray_T6 T6 (
    .CLK(clk),
    .init(init),
    .W0A(T55),
    .W0E(T32),
    .W0I(T24),
    .W0M(T8),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(T5)
  );
  assign T8 = T9;
  assign T9 = {T19, T10};
  assign T10 = {T17, T11};
  assign T11 = 22'h0 - T50;
  assign T50 = {21'h0, T12};
  assign T12 = T13[1'h0];
  assign T13 = rst ? 4'hf : T14;
  assign T14 = io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T51 = reset ? 7'h0 : T15;
  assign T15 = rst ? T16 : rst_cnt;
  assign T16 = rst_cnt + 7'h1;
  assign T17 = 22'h0 - T52;
  assign T52 = {21'h0, T18};
  assign T18 = T13[1'h1];
  assign T19 = {T22, T20};
  assign T20 = 22'h0 - T53;
  assign T53 = {21'h0, T21};
  assign T21 = T13[2'h2];
  assign T22 = 22'h0 - T54;
  assign T54 = {21'h0, T23};
  assign T23 = T13[2'h3];
  assign T24 = T25;
  assign T25 = {T31, T26};
  assign T26 = {wdata, wdata};
  assign wdata = T27;
  assign T27 = {T30, T28};
  assign T28 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T29;
  assign T29 = 2'h0;
  assign T30 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T31 = {wdata, wdata};
  assign T32 = rst | io_write_valid;
  assign T55 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T56;
  assign T56 = {1'h0, io_write_bits_idx};
  assign T34 = io_read_valid ? io_read_bits_idx : R33;
  assign T35 = T5[6'h2b:5'h16];
  assign T36 = {T38, T37};
  assign T37 = T5[7'h41:6'h2c];
  assign T38 = T5[7'h57:7'h42];
  assign io_resp_0_tag = T39;
  assign T39 = T1[5'h15:2'h2];
  assign io_resp_1_coh_state = T40;
  assign T40 = T1[5'h17:5'h16];
  assign io_resp_1_tag = T41;
  assign T41 = T1[6'h2b:5'h18];
  assign io_resp_2_coh_state = T42;
  assign T42 = T1[6'h2d:6'h2c];
  assign io_resp_2_tag = T43;
  assign T43 = T1[7'h41:6'h2e];
  assign io_resp_3_coh_state = T44;
  assign T44 = T1[7'h43:7'h42];
  assign io_resp_3_tag = T45;
  assign T45 = T1[7'h57:7'h44];
  assign io_write_ready = T46;
  assign T46 = rst ^ 1'h1;
  assign io_read_ready = T47;
  assign T47 = T49 & T48;
  assign T48 = io_write_valid ^ 1'h1;
  assign T49 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T16;
    end
    if(io_read_valid) begin
      R33 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    input [3:0] io_in_4_bits_way_en,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    input [3:0] io_in_3_bits_way_en,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    input [3:0] io_in_2_bits_way_en,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[3:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[5:0] T12;
  wire[5:0] T13;
  wire[5:0] T14;
  wire T15;
  wire[5:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_way_en = T3;
  assign T3 = T11 ? io_in_4_bits_way_en : T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T6 = T7[1'h0];
  assign T7 = chosen;
  assign T8 = T9 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T9 = T7[1'h0];
  assign T10 = T7[1'h1];
  assign T11 = T7[2'h2];
  assign io_out_bits_idx = T12;
  assign T12 = T19 ? io_in_4_bits_idx : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T15 = T7[1'h0];
  assign T16 = T17 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T17 = T7[1'h0];
  assign T18 = T7[1'h1];
  assign T19 = T7[2'h2];
  assign io_out_valid = T20;
  assign T20 = T27 ? io_in_4_valid : T21;
  assign T21 = T26 ? T24 : T22;
  assign T22 = T23 ? io_in_1_valid : io_in_0_valid;
  assign T23 = T7[1'h0];
  assign T24 = T25 ? io_in_3_valid : io_in_2_valid;
  assign T25 = T7[1'h0];
  assign T26 = T7[1'h1];
  assign T27 = T7[2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T30;
  assign T30 = T31 & io_out_ready;
  assign T31 = T32 ^ 1'h1;
  assign T32 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T33;
  assign T33 = T34 & io_out_ready;
  assign T34 = T35 ^ 1'h1;
  assign T35 = T36 | io_in_2_valid;
  assign T36 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T40 | io_in_3_valid;
  assign T40 = T41 | io_in_2_valid;
  assign T41 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input [3:0] io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input [3:0] io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_3,
    output[127:0] io_resp_2,
    output[127:0] io_resp_1,
    output[127:0] io_resp_0,
    input  init
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire[127:0] T6;
  wire[63:0] T7;
  wire[127:0] T8;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[7:0] raddr;
  wire[127:0] T10;
  wire[127:0] T11;
  wire[127:0] T12;
  wire[63:0] T13;
  wire[63:0] T140;
  wire T14;
  wire[1:0] T15;
  wire[63:0] T16;
  wire[63:0] T141;
  wire T17;
  wire[127:0] T18;
  wire[127:0] T19;
  wire[63:0] T20;
  wire[63:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[7:0] waddr;
  reg [7:0] R26;
  wire[7:0] T27;
  wire[63:0] T31;
  wire T32;
  wire T33;
  reg [11:0] R34;
  wire[11:0] T35;
  wire[63:0] T36;
  wire[127:0] T37;
  wire[127:0] T38;
  wire[127:0] T39;
  wire[63:0] T40;
  wire[127:0] T41;
  wire T60;
  wire T61;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[63:0] T46;
  wire[63:0] T142;
  wire T47;
  wire[63:0] T48;
  wire[63:0] T143;
  wire T49;
  wire[127:0] T50;
  wire[127:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  reg [7:0] R58;
  wire[7:0] T59;
  wire[63:0] T62;
  wire[127:0] T63;
  wire[127:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire T67;
  wire T68;
  wire[63:0] T69;
  wire[127:0] T70;
  wire[127:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[127:0] T74;
  wire[127:0] T75;
  wire[127:0] T76;
  wire[63:0] T77;
  wire[127:0] T78;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[127:0] T80;
  wire[127:0] T81;
  wire[127:0] T82;
  wire[63:0] T83;
  wire[63:0] T144;
  wire T84;
  wire[1:0] T85;
  wire[63:0] T86;
  wire[63:0] T145;
  wire T87;
  wire[127:0] T88;
  wire[127:0] T89;
  wire[63:0] T90;
  wire[63:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg [7:0] R96;
  wire[7:0] T97;
  wire[63:0] T101;
  wire T102;
  wire T103;
  reg [11:0] R104;
  wire[11:0] T105;
  wire[63:0] T106;
  wire[127:0] T107;
  wire[127:0] T108;
  wire[127:0] T109;
  wire[63:0] T110;
  wire[127:0] T111;
  wire T130;
  wire T131;
  wire[127:0] T113;
  wire[127:0] T114;
  wire[127:0] T115;
  wire[63:0] T116;
  wire[63:0] T146;
  wire T117;
  wire[63:0] T118;
  wire[63:0] T147;
  wire T119;
  wire[127:0] T120;
  wire[127:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  reg [7:0] R128;
  wire[7:0] T129;
  wire[63:0] T132;
  wire[127:0] T133;
  wire[127:0] T134;
  wire[63:0] T135;
  wire[63:0] T136;
  wire T137;
  wire T138;
  wire[63:0] T139;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R26 = {1{$random}};
    R34 = {1{$random}};
    R58 = {1{$random}};
    R96 = {1{$random}};
    R104 = {1{$random}};
    R128 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T36, T2};
  assign T2 = T32 ? T36 : T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = {T31, T7};
  assign T7 = T8[6'h3f:1'h0];
  assign T28 = T29 & io_read_valid;
  assign T29 = T30 != 2'h0;
  assign T30 = io_read_bits_way_en[1'h1:1'h0];
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T9 T9 (
    .CLK(clk),
    .init(init),
    .W0A(waddr),
    .W0E(T22),
    .W0I(T18),
    .W0M(T11),
    .R1A(raddr),
    .R1E(T28),
    .R1O(T8)
  );
  assign T11 = T12;
  assign T12 = {T16, T13};
  assign T13 = 64'h0 - T140;
  assign T140 = {63'h0, T14};
  assign T14 = T15[1'h0];
  assign T15 = io_write_bits_way_en[1'h1:1'h0];
  assign T16 = 64'h0 - T141;
  assign T141 = {63'h0, T17};
  assign T17 = T15[1'h1];
  assign T18 = T19;
  assign T19 = {T21, T20};
  assign T20 = io_write_bits_data[6'h3f:1'h0];
  assign T21 = io_write_bits_data[6'h3f:1'h0];
  assign T22 = T24 & T23;
  assign T23 = io_write_bits_wmask[1'h0];
  assign T24 = T25 & io_write_valid;
  assign T25 = T15 != 2'h0;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T27 = T28 ? raddr : R26;
  assign T31 = T8[7'h7f:7'h40];
  assign T32 = T33;
  assign T33 = R34[2'h3];
  assign T35 = io_read_valid ? io_read_bits_addr : R34;
  assign T36 = T37[6'h3f:1'h0];
  assign T37 = T38;
  assign T38 = T39;
  assign T39 = {T62, T40};
  assign T40 = T41[6'h3f:1'h0];
  assign T60 = T61 & io_read_valid;
  assign T61 = T30 != 2'h0;
  DataArray_T9 T42 (
    .CLK(clk),
    .init(init),
    .W0A(waddr),
    .W0E(T54),
    .W0I(T50),
    .W0M(T44),
    .R1A(raddr),
    .R1E(T60),
    .R1O(T41)
  );
  assign T44 = T45;
  assign T45 = {T48, T46};
  assign T46 = 64'h0 - T142;
  assign T142 = {63'h0, T47};
  assign T47 = T15[1'h0];
  assign T48 = 64'h0 - T143;
  assign T143 = {63'h0, T49};
  assign T49 = T15[1'h1];
  assign T50 = T51;
  assign T51 = {T53, T52};
  assign T52 = io_write_bits_data[7'h7f:7'h40];
  assign T53 = io_write_bits_data[7'h7f:7'h40];
  assign T54 = T56 & T55;
  assign T55 = io_write_bits_wmask[1'h1];
  assign T56 = T57 & io_write_valid;
  assign T57 = T15 != 2'h0;
  assign T59 = T60 ? raddr : R58;
  assign T62 = T41[7'h7f:7'h40];
  assign io_resp_1 = T63;
  assign T63 = T64;
  assign T64 = {T69, T65};
  assign T65 = T67 ? T69 : T66;
  assign T66 = T4[7'h7f:7'h40];
  assign T67 = T68;
  assign T68 = R34[2'h3];
  assign T69 = T37[7'h7f:7'h40];
  assign io_resp_2 = T70;
  assign T70 = T71;
  assign T71 = {T106, T72};
  assign T72 = T102 ? T106 : T73;
  assign T73 = T74[6'h3f:1'h0];
  assign T74 = T75;
  assign T75 = T76;
  assign T76 = {T101, T77};
  assign T77 = T78[6'h3f:1'h0];
  assign T98 = T99 & io_read_valid;
  assign T99 = T100 != 2'h0;
  assign T100 = io_read_bits_way_en[2'h3:2'h2];
  DataArray_T9 T79 (
    .CLK(clk),
    .init(init),
    .W0A(waddr),
    .W0E(T92),
    .W0I(T88),
    .W0M(T81),
    .R1A(raddr),
    .R1E(T98),
    .R1O(T78)
  );
  assign T81 = T82;
  assign T82 = {T86, T83};
  assign T83 = 64'h0 - T144;
  assign T144 = {63'h0, T84};
  assign T84 = T85[1'h0];
  assign T85 = io_write_bits_way_en[2'h3:2'h2];
  assign T86 = 64'h0 - T145;
  assign T145 = {63'h0, T87};
  assign T87 = T85[1'h1];
  assign T88 = T89;
  assign T89 = {T91, T90};
  assign T90 = io_write_bits_data[6'h3f:1'h0];
  assign T91 = io_write_bits_data[6'h3f:1'h0];
  assign T92 = T94 & T93;
  assign T93 = io_write_bits_wmask[1'h0];
  assign T94 = T95 & io_write_valid;
  assign T95 = T85 != 2'h0;
  assign T97 = T98 ? raddr : R96;
  assign T101 = T78[7'h7f:7'h40];
  assign T102 = T103;
  assign T103 = R104[2'h3];
  assign T105 = io_read_valid ? io_read_bits_addr : R104;
  assign T106 = T107[6'h3f:1'h0];
  assign T107 = T108;
  assign T108 = T109;
  assign T109 = {T132, T110};
  assign T110 = T111[6'h3f:1'h0];
  assign T130 = T131 & io_read_valid;
  assign T131 = T100 != 2'h0;
  DataArray_T9 T112 (
    .CLK(clk),
    .init(init),
    .W0A(waddr),
    .W0E(T124),
    .W0I(T120),
    .W0M(T114),
    .R1A(raddr),
    .R1E(T130),
    .R1O(T111)
  );
  assign T114 = T115;
  assign T115 = {T118, T116};
  assign T116 = 64'h0 - T146;
  assign T146 = {63'h0, T117};
  assign T117 = T85[1'h0];
  assign T118 = 64'h0 - T147;
  assign T147 = {63'h0, T119};
  assign T119 = T85[1'h1];
  assign T120 = T121;
  assign T121 = {T123, T122};
  assign T122 = io_write_bits_data[7'h7f:7'h40];
  assign T123 = io_write_bits_data[7'h7f:7'h40];
  assign T124 = T126 & T125;
  assign T125 = io_write_bits_wmask[1'h1];
  assign T126 = T127 & io_write_valid;
  assign T127 = T85 != 2'h0;
  assign T129 = T130 ? raddr : R128;
  assign T132 = T111[7'h7f:7'h40];
  assign io_resp_3 = T133;
  assign T133 = T134;
  assign T134 = {T139, T135};
  assign T135 = T137 ? T139 : T136;
  assign T136 = T74[7'h7f:7'h40];
  assign T137 = T138;
  assign T138 = R104[2'h3];
  assign T139 = T107[7'h7f:7'h40];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T28) begin
      R26 <= raddr;
    end
    if(io_read_valid) begin
      R34 <= io_read_bits_addr;
    end
    if(T60) begin
      R58 <= raddr;
    end
    if(T98) begin
      R96 <= raddr;
    end
    if(io_read_valid) begin
      R104 <= io_read_bits_addr;
    end
    if(T130) begin
      R128 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input [3:0] io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [3:0] io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[11:0] T2;
  wire[11:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[11:0] T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 2'h0 : T0;
  assign T0 = io_in_1_valid ? 2'h1 : T1;
  assign T1 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T4 = T5[1'h0];
  assign T5 = chosen;
  assign T6 = T7 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T7 = T5[1'h0];
  assign T8 = T5[1'h1];
  assign io_out_bits_way_en = T9;
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T11 = T5[1'h0];
  assign T12 = T13 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T13 = T5[1'h0];
  assign T14 = T5[1'h1];
  assign io_out_valid = T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T5[1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T5[1'h0];
  assign T20 = T5[1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_2_valid;
  assign T29 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[127:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[11:0] T3;
  wire[3:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_wmask = T2;
  assign T2 = T1 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T3;
  assign T3 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T4;
  assign T4 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [4:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] wmask;
  wire[63:0] T3;
  wire[31:0] T4;
  wire[15:0] T5;
  wire[7:0] T6;
  wire[7:0] T119;
  wire T7;
  wire[7:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire T28;
  wire[3:0] T29;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T120;
  wire T32;
  wire[15:0] T33;
  wire[7:0] T34;
  wire[7:0] T121;
  wire T35;
  wire[7:0] T36;
  wire[7:0] T122;
  wire T37;
  wire[31:0] T38;
  wire[15:0] T39;
  wire[7:0] T40;
  wire[7:0] T123;
  wire T41;
  wire[7:0] T42;
  wire[7:0] T124;
  wire T43;
  wire[15:0] T44;
  wire[7:0] T45;
  wire[7:0] T125;
  wire T46;
  wire[7:0] T47;
  wire[7:0] T126;
  wire T48;
  wire[63:0] T49;
  wire[63:0] out;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] T55;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[31:0] T58;
  wire T59;
  wire[63:0] T60;
  wire[31:0] T61;
  wire[15:0] T62;
  wire T63;
  wire[63:0] T64;
  wire[31:0] T65;
  wire[15:0] T66;
  wire[7:0] T67;
  wire T68;
  wire T69;
  wire max;
  wire T70;
  wire T71;
  wire min;
  wire T72;
  wire T73;
  wire less;
  wire T74;
  wire cmp_rhs;
  wire T75;
  wire[63:0] rhs;
  wire[63:0] T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire word;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire cmp_lhs;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire sgned;
  wire T94;
  wire T95;
  wire lt;
  wire T96;
  wire T97;
  wire lt_lo;
  wire[31:0] T98;
  wire[31:0] T99;
  wire eq_hi;
  wire[31:0] T100;
  wire[31:0] T101;
  wire lt_hi;
  wire[31:0] T102;
  wire[31:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire[63:0] T107;
  wire T108;
  wire[63:0] T109;
  wire T110;
  wire[63:0] T111;
  wire T112;
  wire[63:0] adder_out;
  wire[63:0] T113;
  wire[63:0] mask;
  wire[63:0] T127;
  wire[31:0] T114;
  wire T115;
  wire[63:0] T116;
  wire[63:0] T117;
  wire T118;


  assign io_out = T0;
  assign T0 = T49 | T1;
  assign T1 = T2 & io_lhs;
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T38, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = 8'h0 - T119;
  assign T119 = {7'h0, T7};
  assign T7 = T8[1'h0];
  assign T8 = {T26, T9};
  assign T9 = T25 ? 4'h0 : T10;
  assign T10 = {T20, T11};
  assign T11 = T19 ? 2'h0 : T12;
  assign T12 = {T15, T13};
  assign T13 = T14 == 1'h0;
  assign T14 = io_addr[1'h0];
  assign T15 = T18 | T16;
  assign T16 = 2'h1 <= T17;
  assign T17 = io_typ[1'h1:1'h0];
  assign T18 = io_addr[1'h0];
  assign T19 = io_addr[1'h1];
  assign T20 = T23 | T21;
  assign T21 = T22 ? 2'h3 : 2'h0;
  assign T22 = 2'h2 <= T17;
  assign T23 = T24 ? T12 : 2'h0;
  assign T24 = io_addr[1'h1];
  assign T25 = io_addr[2'h2];
  assign T26 = T29 | T27;
  assign T27 = T28 ? 4'hf : 4'h0;
  assign T28 = 2'h3 <= T17;
  assign T29 = T30 ? T10 : 4'h0;
  assign T30 = io_addr[2'h2];
  assign T31 = 8'h0 - T120;
  assign T120 = {7'h0, T32};
  assign T32 = T8[1'h1];
  assign T33 = {T36, T34};
  assign T34 = 8'h0 - T121;
  assign T121 = {7'h0, T35};
  assign T35 = T8[2'h2];
  assign T36 = 8'h0 - T122;
  assign T122 = {7'h0, T37};
  assign T37 = T8[2'h3];
  assign T38 = {T44, T39};
  assign T39 = {T42, T40};
  assign T40 = 8'h0 - T123;
  assign T123 = {7'h0, T41};
  assign T41 = T8[3'h4];
  assign T42 = 8'h0 - T124;
  assign T124 = {7'h0, T43};
  assign T43 = T8[3'h5];
  assign T44 = {T47, T45};
  assign T45 = 8'h0 - T125;
  assign T125 = {7'h0, T46};
  assign T46 = T8[3'h6];
  assign T47 = 8'h0 - T126;
  assign T126 = {7'h0, T48};
  assign T48 = T8[3'h7];
  assign T49 = wmask & out;
  assign out = T118 ? adder_out : T50;
  assign T50 = T112 ? T111 : T51;
  assign T51 = T110 ? T109 : T52;
  assign T52 = T108 ? T107 : T53;
  assign T53 = T69 ? io_lhs : T54;
  assign T54 = T68 ? T64 : T55;
  assign T55 = T63 ? T60 : T56;
  assign T56 = T59 ? T57 : io_rhs;
  assign T57 = {T58, T58};
  assign T58 = io_rhs[5'h1f:1'h0];
  assign T59 = T17 == 2'h2;
  assign T60 = {T61, T61};
  assign T61 = {T62, T62};
  assign T62 = io_rhs[4'hf:1'h0];
  assign T63 = T17 == 2'h1;
  assign T64 = {T65, T65};
  assign T65 = {T66, T66};
  assign T66 = {T67, T67};
  assign T67 = io_rhs[3'h7:1'h0];
  assign T68 = T17 == 2'h0;
  assign T69 = less ? min : max;
  assign max = T71 | T70;
  assign T70 = io_cmd == 5'hf;
  assign T71 = io_cmd == 5'hd;
  assign min = T73 | T72;
  assign T72 = io_cmd == 5'he;
  assign T73 = io_cmd == 5'hc;
  assign less = T106 ? lt : T74;
  assign T74 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T80 ? T79 : T75;
  assign T75 = rhs[6'h3f];
  assign rhs = T78 ? T76 : io_rhs;
  assign T76 = {T77, T77};
  assign T77 = io_rhs[5'h1f:1'h0];
  assign T78 = T17 == 2'h2;
  assign T79 = rhs[5'h1f];
  assign T80 = word & T81;
  assign T81 = T82 ^ 1'h1;
  assign T82 = io_addr[2'h2];
  assign word = T84 | T83;
  assign T83 = io_typ == 3'h4;
  assign T84 = T86 | T85;
  assign T85 = io_typ == 3'h0;
  assign T86 = T88 | T87;
  assign T87 = io_typ == 3'h6;
  assign T88 = io_typ == 3'h2;
  assign cmp_lhs = T91 ? T90 : T89;
  assign T89 = io_lhs[6'h3f];
  assign T90 = io_lhs[5'h1f];
  assign T91 = word & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = io_addr[2'h2];
  assign sgned = T95 | T94;
  assign T94 = io_cmd == 5'hd;
  assign T95 = io_cmd == 5'hc;
  assign lt = word ? T104 : T96;
  assign T96 = lt_hi | T97;
  assign T97 = eq_hi & lt_lo;
  assign lt_lo = T99 < T98;
  assign T98 = rhs[5'h1f:1'h0];
  assign T99 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T101 == T100;
  assign T100 = rhs[6'h3f:6'h20];
  assign T101 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T103 < T102;
  assign T102 = rhs[6'h3f:6'h20];
  assign T103 = io_lhs[6'h3f:6'h20];
  assign T104 = T105 ? lt_hi : lt_lo;
  assign T105 = io_addr[2'h2];
  assign T106 = cmp_lhs == cmp_rhs;
  assign T107 = io_lhs ^ rhs;
  assign T108 = io_cmd == 5'h9;
  assign T109 = io_lhs | rhs;
  assign T110 = io_cmd == 5'ha;
  assign T111 = io_lhs & rhs;
  assign T112 = io_cmd == 5'hb;
  assign adder_out = T116 + T113;
  assign T113 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T127;
  assign T127 = {32'h0, T114};
  assign T114 = T115 << 5'h1f;
  assign T115 = io_addr[2'h2];
  assign T116 = T117;
  assign T117 = io_lhs & mask;
  assign T118 = io_cmd == 5'h8;
endmodule

module LockingArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [5:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_voluntary,
    input [2:0] io_in_1_bits_r_type,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [5:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_voluntary,
    input [2:0] io_in_0_bits_r_type,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[5:0] io_out_bits_client_xact_id,
    output io_out_bits_voluntary,
    output[2:0] io_out_bits_r_type,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T37;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T38;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T39;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire[127:0] T22;
  wire T23;
  wire[2:0] T24;
  wire T25;
  wire[5:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T37 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T12 & T7;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_out_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_out_bits_r_type;
  assign T11 = 3'h0 == io_out_bits_r_type;
  assign T12 = io_out_valid & io_out_ready;
  assign T38 = reset ? 1'h0 : T13;
  assign T13 = T20 ? 1'h0 : T14;
  assign T14 = T6 ? T15 : locked;
  assign T15 = T16 ^ 1'h1;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T39 = reset ? 2'h0 : T19;
  assign T19 = T6 ? T17 : R18;
  assign T20 = T12 & T21;
  assign T21 = T7 ^ 1'h1;
  assign io_out_bits_data = T22;
  assign T22 = T23 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T23 = chosen;
  assign io_out_bits_r_type = T24;
  assign T24 = T23 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_voluntary = T25;
  assign T25 = T23 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_client_xact_id = T26;
  assign T26 = T23 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T27;
  assign T27 = T23 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T28;
  assign T28 = T23 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T29;
  assign T29 = T23 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T30;
  assign T30 = T31 & io_out_ready;
  assign T31 = locked ? T32 : 1'h1;
  assign T32 = lockIdx == 1'h0;
  assign io_in_1_ready = T33;
  assign T33 = T34 & io_out_ready;
  assign T34 = locked ? T36 : T35;
  assign T35 = io_in_0_valid ^ 1'h1;
  assign T36 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T20) begin
      locked <= 1'h0;
    end else if(T6) begin
      locked <= T15;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T6) begin
      R18 <= T17;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_addr,
    input [9:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_kill,
    input  io_cpu_req_bits_phys,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_addr,
    output[9:0] io_cpu_resp_bits_tag,
    output[4:0] io_cpu_resp_bits_cmd,
    output[2:0] io_cpu_resp_bits_typ,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_word_bypass,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[9:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_invalidate_lr,
    output io_cpu_ordered,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[5:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [5:0] io_mem_grant_bits_client_xact_id,
    input [3:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [25:0] io_mem_probe_bits_addr_block,
    input [1:0] io_mem_probe_bits_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_addr_beat,
    output[25:0] io_mem_release_bits_addr_block,
    output[5:0] io_mem_release_bits_client_xact_id,
    output io_mem_release_bits_voluntary,
    output[2:0] io_mem_release_bits_r_type,
    output[127:0] io_mem_release_bits_data,
    input  init
);

  reg  T0;
  wire T1;
  wire T2;
  wire T3;
  reg  R4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg [63:0] s2_req_data;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  s1_replay;
  wire T559;
  wire T20;
  wire T21;
  wire s1_write;
  wire T22;
  wire T23;
  reg [4:0] s1_req_cmd;
  wire[4:0] T24;
  wire[4:0] T25;
  wire[4:0] T26;
  reg [4:0] s2_req_cmd;
  wire[4:0] T27;
  wire s2_recycle;
  wire T28;
  reg  s2_recycle_next;
  wire T560;
  wire T29;
  wire T30;
  reg  s1_valid;
  wire T561;
  wire T31;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire[1:0] T32;
  wire T33;
  wire s2_hit;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  reg [1:0] R48;
  wire[1:0] T49;
  wire T50;
  reg [3:0] s2_tag_match_way;
  wire[3:0] T51;
  wire[3:0] s1_tag_match_way;
  wire[3:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[3:0] s1_tag_eq_way;
  wire[3:0] T57;
  wire[1:0] T58;
  wire T59;
  wire[19:0] T60;
  wire[31:0] s1_addr;
  wire[11:0] T61;
  reg [39:0] s1_req_addr;
  wire[39:0] T62;
  wire[39:0] T63;
  wire[39:0] T64;
  wire[39:0] T65;
  wire[39:0] T66;
  wire[39:0] T562;
  wire[31:0] T67;
  wire[25:0] T68;
  wire[39:0] T563;
  wire[31:0] T69;
  wire[25:0] T70;
  reg [39:0] s2_req_addr;
  wire[39:0] T71;
  wire[39:0] T564;
  wire T72;
  wire[19:0] T73;
  wire[1:0] T74;
  wire T75;
  wire[19:0] T76;
  wire T77;
  wire[19:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  reg [1:0] R92;
  wire[1:0] T93;
  wire T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  reg [1:0] R98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T101;
  wire[1:0] T102;
  reg [1:0] R103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire s2_tag_match;
  wire T127;
  wire s2_replay;
  wire T128;
  reg  R129;
  wire T565;
  reg  s2_valid;
  wire T566;
  wire s1_valid_masked;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire T138;
  reg  s1_recycled;
  wire T567;
  wire T139;
  wire[63:0] T568;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T140;
  wire[63:0] T141;
  wire[127:0] s2_data_muxed;
  wire[127:0] T142;
  wire[127:0] s2_data_3;
  wire[127:0] T143;
  wire[127:0] T144;
  reg [63:0] R145;
  wire[63:0] T569;
  wire[127:0] T146;
  wire[127:0] T570;
  wire[127:0] T147;
  wire T148;
  wire T149;
  reg [63:0] R150;
  wire[63:0] T151;
  wire[63:0] T152;
  wire T153;
  wire s1_writeback;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire[127:0] T158;
  wire[127:0] T159;
  wire[127:0] s2_data_2;
  wire[127:0] T160;
  wire[127:0] T161;
  reg [63:0] R162;
  wire[63:0] T571;
  wire[127:0] T163;
  wire[127:0] T572;
  wire[127:0] T164;
  wire T165;
  wire T166;
  reg [63:0] R167;
  wire[63:0] T168;
  wire[63:0] T169;
  wire T170;
  wire T171;
  wire[127:0] T172;
  wire[127:0] T173;
  wire[127:0] s2_data_1;
  wire[127:0] T174;
  wire[127:0] T175;
  reg [63:0] R176;
  wire[63:0] T573;
  wire[127:0] T177;
  wire[127:0] T574;
  wire[127:0] T178;
  wire T179;
  wire T180;
  reg [63:0] R181;
  wire[63:0] T182;
  wire[63:0] T183;
  wire T184;
  wire T185;
  wire[127:0] T186;
  wire[127:0] s2_data_0;
  wire[127:0] T187;
  wire[127:0] T188;
  reg [63:0] R189;
  wire[63:0] T575;
  wire[127:0] T190;
  wire[127:0] T576;
  wire[127:0] T191;
  wire T192;
  wire T193;
  reg [63:0] R194;
  wire[63:0] T195;
  wire[63:0] T196;
  wire T197;
  wire T198;
  wire[63:0] T199;
  wire[127:0] T577;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  reg [63:0] s4_req_data;
  wire[63:0] T203;
  wire T204;
  reg  s3_valid;
  wire T578;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire s2_sc_fail;
  wire T215;
  wire s2_lrsc_addr_match;
  wire T216;
  wire[33:0] T217;
  reg [33:0] lrsc_addr;
  wire[33:0] T218;
  wire[33:0] T219;
  wire T220;
  wire s2_lr;
  wire T221;
  wire T222;
  wire s2_valid_masked;
  wire T223;
  wire T224;
  wire s2_nack;
  wire s2_nack_miss;
  wire T225;
  wire T226;
  wire T227;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T228;
  wire s1_nack;
  wire T229;
  wire T230;
  wire T231;
  wire[5:0] T232;
  wire T233;
  wire T234;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T579;
  wire[4:0] T235;
  wire[4:0] T236;
  wire[4:0] T237;
  wire[4:0] T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire s2_sc;
  wire T243;
  wire T244;
  reg [63:0] s3_req_data;
  wire[63:0] T580;
  wire[127:0] T245;
  wire[127:0] T581;
  wire[63:0] T246;
  wire[127:0] T247;
  wire[127:0] T582;
  wire[127:0] s2_data_corrected;
  wire[127:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  reg [4:0] s3_req_cmd;
  wire[4:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[36:0] T270;
  reg [39:0] s3_req_addr;
  wire[39:0] T271;
  wire[36:0] T583;
  wire[28:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire[36:0] T283;
  wire[36:0] T584;
  wire[28:0] T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  reg [4:0] s4_req_cmd;
  wire[4:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[36:0] T301;
  reg [39:0] s4_req_addr;
  wire[39:0] T302;
  wire[36:0] T585;
  wire[28:0] T303;
  reg  s4_valid;
  wire T586;
  wire T304;
  reg  s2_store_bypass;
  wire T305;
  wire T306;
  reg [2:0] s2_req_typ;
  wire[2:0] T307;
  reg [2:0] s1_req_typ;
  wire[2:0] T308;
  wire[2:0] T309;
  wire[2:0] T310;
  wire[5:0] T587;
  wire[127:0] T311;
  wire[1:0] rowWMask;
  wire rowIdx;
  wire T312;
  wire[11:0] T588;
  reg [3:0] s3_way;
  wire[3:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire[11:0] T589;
  wire[11:0] T590;
  wire[11:0] T591;
  wire[127:0] T326;
  wire[127:0] T327;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[5:0] T592;
  wire[33:0] T328;
  wire[5:0] T593;
  wire[33:0] T329;
  reg  s1_req_phys;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  reg  s2_req_phys;
  wire T335;
  wire[27:0] T336;
  wire T337;
  wire T338;
  wire T339;
  wire s1_readwrite;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire s1_read;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire cache_pass;
  wire T354;
  reg  s2_killed;
  wire T355;
  wire[3:0] T356;
  wire[3:0] s2_replaced_way_en;
  reg [1:0] R357;
  wire[1:0] T358;
  wire[1:0] T359;
  reg [15:0] R360;
  wire[15:0] T594;
  wire[15:0] T361;
  wire[15:0] T362;
  wire[14:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire[1:0] T373;
  wire[1:0] T374;
  wire[21:0] T375;
  wire[21:0] T376;
  wire[21:0] T377;
  wire[21:0] T378;
  reg [1:0] R379;
  wire[1:0] T380;
  wire T381;
  wire T382;
  wire[3:0] s1_replaced_way_en;
  wire[1:0] T383;
  reg [19:0] R384;
  wire[19:0] T385;
  wire T386;
  wire[21:0] T387;
  wire[21:0] T388;
  wire[21:0] T389;
  wire[21:0] T390;
  reg [1:0] R391;
  wire[1:0] T392;
  wire T393;
  wire T394;
  reg [19:0] R395;
  wire[19:0] T396;
  wire T397;
  wire[21:0] T398;
  wire[21:0] T399;
  wire[21:0] T400;
  wire[21:0] T401;
  reg [1:0] R402;
  wire[1:0] T403;
  wire T404;
  wire T405;
  reg [19:0] R406;
  wire[19:0] T407;
  wire T408;
  wire[21:0] T409;
  wire[21:0] T410;
  wire[21:0] T411;
  reg [1:0] R412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  reg [19:0] R416;
  wire[19:0] T417;
  wire T418;
  wire[1:0] T419;
  wire[19:0] T420;
  wire[19:0] T421;
  wire[19:0] T422;
  reg  s2_req_kill;
  wire T423;
  reg  s1_req_kill;
  wire T424;
  wire T425;
  wire T426;
  reg [9:0] s2_req_tag;
  wire[9:0] T427;
  reg [9:0] s1_req_tag;
  wire[9:0] T428;
  wire[9:0] T429;
  wire[9:0] T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire misaligned;
  wire[39:0] T467;
  wire[39:0] T595;
  wire[2:0] T468;
  wire[3:0] T469;
  wire[3:0] T470;
  wire[1:0] T471;
  wire T472;
  wire T473;
  wire[63:0] T474;
  wire[63:0] uncache_resp_bits_store_data;
  wire[63:0] cache_resp_bits_store_data;
  wire[63:0] T475;
  wire[31:0] T476;
  wire[31:0] T477;
  wire[31:0] T478;
  wire T479;
  wire[31:0] T480;
  wire[31:0] T481;
  wire[31:0] T482;
  wire[31:0] T596;
  wire T483;
  wire T484;
  wire T485;
  wire[2:0] T486;
  wire T487;
  wire[1:0] T488;
  wire T489;
  wire uncache_resp_bits_has_data;
  wire cache_resp_bits_has_data;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire uncache_resp_bits_replay;
  wire cache_resp_bits_replay;
  wire T500;
  wire uncache_resp_bits_nack;
  wire cache_resp_bits_nack;
  wire T501;
  wire[63:0] T502;
  wire[63:0] uncache_resp_bits_data;
  wire[63:0] cache_resp_bits_data;
  wire[63:0] T503;
  wire[63:0] T597;
  wire[63:0] T504;
  wire[7:0] T505;
  wire[7:0] T506;
  wire[7:0] T507;
  wire[63:0] T508;
  wire[15:0] T509;
  wire[15:0] T510;
  wire[63:0] T511;
  wire[31:0] T512;
  wire[31:0] T513;
  wire[31:0] T514;
  wire T515;
  wire[31:0] T516;
  wire[31:0] T517;
  wire[31:0] T518;
  wire[31:0] T598;
  wire T519;
  wire T520;
  wire T521;
  wire[15:0] T522;
  wire T523;
  wire[47:0] T524;
  wire[47:0] T525;
  wire[47:0] T526;
  wire[47:0] T599;
  wire T527;
  wire T528;
  wire T529;
  wire[7:0] T530;
  wire T531;
  wire[55:0] T532;
  wire[55:0] T533;
  wire[55:0] T534;
  wire[55:0] T600;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire[2:0] T539;
  wire[2:0] uncache_resp_bits_typ;
  wire[2:0] cache_resp_bits_typ;
  wire[4:0] T540;
  wire[4:0] uncache_resp_bits_cmd;
  wire[4:0] cache_resp_bits_cmd;
  wire[9:0] T541;
  wire[9:0] uncache_resp_bits_tag;
  wire[9:0] cache_resp_bits_tag;
  wire[39:0] T542;
  wire[39:0] uncache_resp_bits_addr;
  wire[39:0] cache_resp_bits_addr;
  wire T543;
  wire uncache_resp_valid;
  wire cache_resp_valid;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  reg  block_miss;
  wire T601;
  wire T557;
  wire T558;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire[3:0] wb_io_data_req_bits_way_en;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[1:0] wb_io_release_bits_addr_beat;
  wire[25:0] wb_io_release_bits_addr_block;
  wire[5:0] wb_io_release_bits_client_xact_id;
  wire wb_io_release_bits_voluntary;
  wire[2:0] wb_io_release_bits_r_type;
  wire[127:0] wb_io_release_bits_data;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[1:0] prober_io_rep_bits_addr_beat;
  wire[25:0] prober_io_rep_bits_addr_block;
  wire[5:0] prober_io_rep_bits_client_xact_id;
  wire prober_io_rep_bits_voluntary;
  wire[2:0] prober_io_rep_bits_r_type;
  wire[127:0] prober_io_rep_bits_data;
  wire prober_io_meta_read_valid;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire[3:0] prober_io_meta_write_bits_way_en;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[1:0] prober_io_wb_req_bits_addr_beat;
  wire[25:0] prober_io_wb_req_bits_addr_block;
  wire[5:0] prober_io_wb_req_bits_client_xact_id;
  wire prober_io_wb_req_bits_voluntary;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire[127:0] prober_io_wb_req_bits_data;
  wire[3:0] prober_io_wb_req_bits_way_en;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[19:0] meta_io_resp_3_tag;
  wire[1:0] meta_io_resp_3_coh_state;
  wire[19:0] meta_io_resp_2_tag;
  wire[1:0] meta_io_resp_2_coh_state;
  wire[19:0] meta_io_resp_1_tag;
  wire[1:0] meta_io_resp_1_coh_state;
  wire[19:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  wire[3:0] metaReadArb_io_out_bits_way_en;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire[3:0] metaWriteArb_io_out_bits_way_en;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_3;
  wire[127:0] data_io_resp_2;
  wire[127:0] data_io_resp_1;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire[3:0] readArb_io_out_bits_way_en;
  wire[11:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire[3:0] writeArb_io_out_bits_way_en;
  wire[11:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[1:0] releaseArb_io_out_bits_addr_beat;
  wire[25:0] releaseArb_io_out_bits_addr_block;
  wire[5:0] releaseArb_io_out_bits_client_xact_id;
  wire releaseArb_io_out_bits_voluntary;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire[127:0] releaseArb_io_out_bits_data;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[1:0] FlowThroughSerializer_io_out_bits_addr_beat;
  wire[5:0] FlowThroughSerializer_io_out_bits_client_xact_id;
  wire[3:0] FlowThroughSerializer_io_out_bits_manager_xact_id;
  wire FlowThroughSerializer_io_out_bits_is_builtin_type;
  wire[3:0] FlowThroughSerializer_io_out_bits_g_type;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[1:0] wbArb_io_out_bits_addr_beat;
  wire[25:0] wbArb_io_out_bits_addr_block;
  wire[5:0] wbArb_io_out_bits_client_xact_id;
  wire wbArb_io_out_bits_voluntary;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire[127:0] wbArb_io_out_bits_data;
  wire[3:0] wbArb_io_out_bits_way_en;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[19:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[26:0] dtlb_io_ptw_req_bits_addr;
  wire[1:0] dtlb_io_ptw_req_bits_prv;
  wire dtlb_io_ptw_req_bits_store;
  wire dtlb_io_ptw_req_bits_fetch;
  wire mshrs_io_req_ready;
  wire mshrs_io_resp_valid;
  wire[39:0] mshrs_io_resp_bits_addr;
  wire[9:0] mshrs_io_resp_bits_tag;
  wire[4:0] mshrs_io_resp_bits_cmd;
  wire[2:0] mshrs_io_resp_bits_typ;
  wire[63:0] mshrs_io_resp_bits_data;
  wire mshrs_io_resp_bits_nack;
  wire mshrs_io_resp_bits_replay;
  wire mshrs_io_resp_bits_has_data;
  wire[63:0] mshrs_io_resp_bits_store_data;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr_block;
  wire[5:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[1:0] mshrs_io_mem_req_bits_addr_beat;
  wire mshrs_io_mem_req_bits_is_builtin_type;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[16:0] mshrs_io_mem_req_bits_union;
  wire[127:0] mshrs_io_mem_req_bits_data;
  wire[3:0] mshrs_io_refill_way_en;
  wire[11:0] mshrs_io_refill_addr;
  wire mshrs_io_meta_read_valid;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire[3:0] mshrs_io_meta_read_bits_way_en;
  wire mshrs_io_meta_write_valid;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire[3:0] mshrs_io_meta_write_bits_way_en;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire[39:0] mshrs_io_replay_bits_addr;
  wire[9:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_kill;
  wire mshrs_io_replay_bits_phys;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_wb_req_valid;
  wire[1:0] mshrs_io_wb_req_bits_addr_beat;
  wire[25:0] mshrs_io_wb_req_bits_addr_block;
  wire[5:0] mshrs_io_wb_req_bits_client_xact_id;
  wire mshrs_io_wb_req_bits_voluntary;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire[127:0] mshrs_io_wb_req_bits_data;
  wire[3:0] mshrs_io_wb_req_bits_way_en;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {1{$random}};
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    R48 = {1{$random}};
    s2_tag_match_way = {1{$random}};
    s1_req_addr = {2{$random}};
    s2_req_addr = {2{$random}};
    R92 = {1{$random}};
    R98 = {1{$random}};
    R103 = {1{$random}};
    R129 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R145 = {2{$random}};
    R150 = {2{$random}};
    R162 = {2{$random}};
    R167 = {2{$random}};
    R176 = {2{$random}};
    R181 = {2{$random}};
    R189 = {2{$random}};
    R194 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    s2_killed = {1{$random}};
    R357 = {1{$random}};
    R360 = {1{$random}};
    R379 = {1{$random}};
    R384 = {1{$random}};
    R391 = {1{$random}};
    R395 = {1{$random}};
    R402 = {1{$random}};
    R406 = {1{$random}};
    R412 = {1{$random}};
    R416 = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    block_miss = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = R4 & io_cpu_resp_valid;
  assign T5 = T6 | io_cpu_xcpt_pf_st;
  assign T6 = T7 | io_cpu_xcpt_pf_ld;
  assign T7 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T8 = writeArb_io_in_1_ready | T9;
  assign T9 = T10 ^ 1'h1;
  assign T10 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T14 : T11;
  assign T11 = T13 | T12;
  assign T12 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T13 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T14 = T16 | T15;
  assign T15 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T16 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T17 = T138 ? s1_req_data : T18;
  assign T18 = T21 ? T19 : s2_req_data;
  assign T19 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T559 = reset ? 1'h0 : T20;
  assign T20 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T21 = s1_clk_en & s1_write;
  assign s1_write = T132 | T22;
  assign T22 = T131 | T23;
  assign T23 = s1_req_cmd == 5'h4;
  assign T24 = s2_recycle ? s2_req_cmd : T25;
  assign T25 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T26;
  assign T26 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T27 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T28;
  assign T28 = s2_recycle_ecc | s2_recycle_next;
  assign T560 = reset ? 1'h0 : T29;
  assign T29 = T30 ? s2_recycle_ecc : s2_recycle_next;
  assign T30 = s1_valid | s1_replay;
  assign T561 = reset ? 1'h0 : T31;
  assign T31 = io_cpu_req_ready & io_cpu_req_valid;
  assign s2_recycle_ecc = T33 & s2_data_correctable;
  assign s2_data_correctable = T32[1'h0];
  assign T32 = 2'h0;
  assign T33 = T127 & s2_hit;
  assign s2_hit = T106 & T34;
  assign T34 = T44 == T35;
  assign T35 = T36;
  assign T36 = T37 ? 2'h3 : T44;
  assign T37 = T41 | T38;
  assign T38 = T40 | T39;
  assign T39 = s2_req_cmd == 5'h4;
  assign T40 = s2_req_cmd[2'h3];
  assign T41 = T43 | T42;
  assign T42 = s2_req_cmd == 5'h7;
  assign T43 = s2_req_cmd == 5'h1;
  assign T44 = T45;
  assign T45 = T89 | T46;
  assign T46 = T50 ? T47 : 2'h0;
  assign T47 = R48;
  assign T49 = s1_clk_en ? meta_io_resp_3_coh_state : R48;
  assign T50 = s2_tag_match_way[2'h3];
  assign T51 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T52;
  assign T52 = {T82, T53};
  assign T53 = {T79, T54};
  assign T54 = T56 & T55;
  assign T55 = meta_io_resp_0_coh_state != 2'h0;
  assign T56 = s1_tag_eq_way[1'h0];
  assign s1_tag_eq_way = T57;
  assign T57 = {T74, T58};
  assign T58 = {T72, T59};
  assign T59 = meta_io_resp_0_tag == T60;
  assign T60 = s1_addr >> 4'hc;
  assign s1_addr = {dtlb_io_resp_ppn, T61};
  assign T61 = s1_req_addr[4'hb:1'h0];
  assign T62 = s2_recycle ? s2_req_addr : T63;
  assign T63 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T64;
  assign T64 = prober_io_meta_read_valid ? T563 : T65;
  assign T65 = wb_io_meta_read_valid ? T562 : T66;
  assign T66 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T562 = {8'h0, T67};
  assign T67 = T68 << 3'h6;
  assign T68 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T563 = {8'h0, T69};
  assign T69 = T70 << 3'h6;
  assign T70 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T71 = s1_clk_en ? T564 : s2_req_addr;
  assign T564 = {8'h0, s1_addr};
  assign T72 = meta_io_resp_1_tag == T73;
  assign T73 = s1_addr >> 4'hc;
  assign T74 = {T77, T75};
  assign T75 = meta_io_resp_2_tag == T76;
  assign T76 = s1_addr >> 4'hc;
  assign T77 = meta_io_resp_3_tag == T78;
  assign T78 = s1_addr >> 4'hc;
  assign T79 = T81 & T80;
  assign T80 = meta_io_resp_1_coh_state != 2'h0;
  assign T81 = s1_tag_eq_way[1'h1];
  assign T82 = {T86, T83};
  assign T83 = T85 & T84;
  assign T84 = meta_io_resp_2_coh_state != 2'h0;
  assign T85 = s1_tag_eq_way[2'h2];
  assign T86 = T88 & T87;
  assign T87 = meta_io_resp_3_coh_state != 2'h0;
  assign T88 = s1_tag_eq_way[2'h3];
  assign T89 = T95 | T90;
  assign T90 = T94 ? T91 : 2'h0;
  assign T91 = R92;
  assign T93 = s1_clk_en ? meta_io_resp_2_coh_state : R92;
  assign T94 = s2_tag_match_way[2'h2];
  assign T95 = T101 | T96;
  assign T96 = T100 ? T97 : 2'h0;
  assign T97 = R98;
  assign T99 = s1_clk_en ? meta_io_resp_1_coh_state : R98;
  assign T100 = s2_tag_match_way[1'h1];
  assign T101 = T105 ? T102 : 2'h0;
  assign T102 = R103;
  assign T104 = s1_clk_en ? meta_io_resp_0_coh_state : R103;
  assign T105 = s2_tag_match_way[1'h0];
  assign T106 = s2_tag_match & T107;
  assign T107 = T116 ? T113 : T108;
  assign T108 = T110 | T109;
  assign T109 = 2'h3 == T44;
  assign T110 = T112 | T111;
  assign T111 = 2'h2 == T44;
  assign T112 = 2'h1 == T44;
  assign T113 = T115 | T114;
  assign T114 = 2'h3 == T44;
  assign T115 = 2'h2 == T44;
  assign T116 = T118 | T117;
  assign T117 = s2_req_cmd == 5'h6;
  assign T118 = T120 | T119;
  assign T119 = s2_req_cmd == 5'h3;
  assign T120 = T124 | T121;
  assign T121 = T123 | T122;
  assign T122 = s2_req_cmd == 5'h4;
  assign T123 = s2_req_cmd[2'h3];
  assign T124 = T126 | T125;
  assign T125 = s2_req_cmd == 5'h7;
  assign T126 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign T127 = s2_valid | s2_replay;
  assign s2_replay = R129 & T128;
  assign T128 = s2_req_cmd != 5'h5;
  assign T565 = reset ? 1'h0 : s1_replay;
  assign T566 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T130;
  assign T130 = io_cpu_req_bits_kill ^ 1'h1;
  assign T131 = s1_req_cmd[2'h3];
  assign T132 = T134 | T133;
  assign T133 = s1_req_cmd == 5'h7;
  assign T134 = s1_req_cmd == 5'h1;
  assign T135 = s2_recycle ? s2_req_data : T136;
  assign T136 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T137;
  assign T137 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T138 = s1_clk_en & s1_recycled;
  assign T567 = reset ? 1'h0 : T139;
  assign T139 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T568 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T577 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> 7'h0;
  assign s2_data_uncorrected = T140;
  assign T140 = {T199, T141};
  assign T141 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T158 | T142;
  assign T142 = T157 ? s2_data_3 : 128'h0;
  assign s2_data_3 = T143;
  assign T143 = T144;
  assign T144 = {R150, R145};
  assign T569 = T146[6'h3f:1'h0];
  assign T146 = T148 ? T147 : T570;
  assign T570 = {64'h0, R145};
  assign T147 = data_io_resp_3 >> 1'h0;
  assign T148 = s1_clk_en & T149;
  assign T149 = s1_tag_eq_way[2'h3];
  assign T151 = T153 ? T152 : R150;
  assign T152 = data_io_resp_3 >> 7'h40;
  assign T153 = T148 & s1_writeback;
  assign s1_writeback = T155 & T154;
  assign T154 = s1_replay ^ 1'h1;
  assign T155 = s1_clk_en & T156;
  assign T156 = s1_valid ^ 1'h1;
  assign T157 = s2_tag_match_way[2'h3];
  assign T158 = T172 | T159;
  assign T159 = T171 ? s2_data_2 : 128'h0;
  assign s2_data_2 = T160;
  assign T160 = T161;
  assign T161 = {R167, R162};
  assign T571 = T163[6'h3f:1'h0];
  assign T163 = T165 ? T164 : T572;
  assign T572 = {64'h0, R162};
  assign T164 = data_io_resp_2 >> 1'h0;
  assign T165 = s1_clk_en & T166;
  assign T166 = s1_tag_eq_way[2'h2];
  assign T168 = T170 ? T169 : R167;
  assign T169 = data_io_resp_2 >> 7'h40;
  assign T170 = T165 & s1_writeback;
  assign T171 = s2_tag_match_way[2'h2];
  assign T172 = T186 | T173;
  assign T173 = T185 ? s2_data_1 : 128'h0;
  assign s2_data_1 = T174;
  assign T174 = T175;
  assign T175 = {R181, R176};
  assign T573 = T177[6'h3f:1'h0];
  assign T177 = T179 ? T178 : T574;
  assign T574 = {64'h0, R176};
  assign T178 = data_io_resp_1 >> 1'h0;
  assign T179 = s1_clk_en & T180;
  assign T180 = s1_tag_eq_way[1'h1];
  assign T182 = T184 ? T183 : R181;
  assign T183 = data_io_resp_1 >> 7'h40;
  assign T184 = T179 & s1_writeback;
  assign T185 = s2_tag_match_way[1'h1];
  assign T186 = T198 ? s2_data_0 : 128'h0;
  assign s2_data_0 = T187;
  assign T187 = T188;
  assign T188 = {R194, R189};
  assign T575 = T190[6'h3f:1'h0];
  assign T190 = T192 ? T191 : T576;
  assign T576 = {64'h0, R189};
  assign T191 = data_io_resp_0 >> 1'h0;
  assign T192 = s1_clk_en & T193;
  assign T193 = s1_tag_eq_way[1'h0];
  assign T195 = T197 ? T196 : R194;
  assign T196 = data_io_resp_0 >> 7'h40;
  assign T197 = T192 & s1_writeback;
  assign T198 = s2_tag_match_way[1'h0];
  assign T199 = s2_data_muxed[7'h7f:7'h40];
  assign T577 = {64'h0, s2_store_bypass_data};
  assign T200 = T288 ? T201 : s2_store_bypass_data;
  assign T201 = T273 ? amoalu_io_out : T202;
  assign T202 = T259 ? s3_req_data : s4_req_data;
  assign T203 = T204 ? s3_req_data : s4_req_data;
  assign T204 = s3_valid & metaReadArb_io_out_valid;
  assign T578 = reset ? 1'h0 : T205;
  assign T205 = T213 & T206;
  assign T206 = T210 | T207;
  assign T207 = T209 | T208;
  assign T208 = s2_req_cmd == 5'h4;
  assign T209 = s2_req_cmd[2'h3];
  assign T210 = T212 | T211;
  assign T211 = s2_req_cmd == 5'h7;
  assign T212 = s2_req_cmd == 5'h1;
  assign T213 = T243 & T214;
  assign T214 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T215;
  assign T215 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T216;
  assign T216 = lrsc_addr == T217;
  assign T217 = s2_req_addr >> 3'h6;
  assign T218 = T220 ? T219 : lrsc_addr;
  assign T219 = s2_req_addr >> 3'h6;
  assign T220 = T221 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T221 = T222 | s2_replay;
  assign T222 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T223;
  assign T223 = s2_valid & T224;
  assign T224 = s2_nack ^ 1'h1;
  assign s2_nack = T227 | s2_nack_miss;
  assign s2_nack_miss = T226 & T225;
  assign T225 = mshrs_io_req_ready ^ 1'h1;
  assign T226 = s2_hit ^ 1'h1;
  assign T227 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T228 = T234 ? s1_nack : s2_nack_hit;
  assign s1_nack = T233 | T229;
  assign T229 = T231 & T230;
  assign T230 = prober_io_req_ready ^ 1'h1;
  assign T231 = T232 == prober_io_meta_write_bits_idx;
  assign T232 = s1_req_addr[4'hb:3'h6];
  assign T233 = T337 & dtlb_io_resp_miss;
  assign T234 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T579 = reset ? 5'h0 : T235;
  assign T235 = io_cpu_invalidate_lr ? 5'h0 : T236;
  assign T236 = T242 ? 5'h0 : T237;
  assign T237 = T240 ? 5'h1f : T238;
  assign T238 = lrsc_valid ? T239 : lrsc_count;
  assign T239 = lrsc_count - 5'h1;
  assign T240 = T220 & T241;
  assign T241 = lrsc_valid ^ 1'h1;
  assign T242 = T221 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T243 = T244 | s2_replay;
  assign T244 = s2_valid_masked & s2_hit;
  assign T580 = T245[6'h3f:1'h0];
  assign T245 = T249 ? T247 : T581;
  assign T581 = {64'h0, T246};
  assign T246 = T249 ? s2_req_data : s3_req_data;
  assign T247 = s2_data_correctable ? s2_data_corrected : T582;
  assign T582 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T248;
  assign T248 = {T199, T141};
  assign T249 = T258 & T250;
  assign T250 = T251 | s2_data_correctable;
  assign T251 = T255 | T252;
  assign T252 = T254 | T253;
  assign T253 = s2_req_cmd == 5'h4;
  assign T254 = s2_req_cmd[2'h3];
  assign T255 = T257 | T256;
  assign T256 = s2_req_cmd == 5'h7;
  assign T257 = s2_req_cmd == 5'h1;
  assign T258 = s2_valid | s2_replay;
  assign T259 = T268 & T260;
  assign T260 = T265 | T261;
  assign T261 = T264 | T262;
  assign T262 = s3_req_cmd == 5'h4;
  assign T263 = T249 ? s2_req_cmd : s3_req_cmd;
  assign T264 = s3_req_cmd[2'h3];
  assign T265 = T267 | T266;
  assign T266 = s3_req_cmd == 5'h7;
  assign T267 = s3_req_cmd == 5'h1;
  assign T268 = s3_valid & T269;
  assign T269 = T583 == T270;
  assign T270 = s3_req_addr >> 2'h3;
  assign T271 = T249 ? s2_req_addr : s3_req_addr;
  assign T583 = {8'h0, T272};
  assign T272 = s1_addr >> 2'h3;
  assign T273 = T281 & T274;
  assign T274 = T278 | T275;
  assign T275 = T277 | T276;
  assign T276 = s2_req_cmd == 5'h4;
  assign T277 = s2_req_cmd[2'h3];
  assign T278 = T280 | T279;
  assign T279 = s2_req_cmd == 5'h7;
  assign T280 = s2_req_cmd == 5'h1;
  assign T281 = T285 & T282;
  assign T282 = T584 == T283;
  assign T283 = s2_req_addr >> 2'h3;
  assign T584 = {8'h0, T284};
  assign T284 = s1_addr >> 2'h3;
  assign T285 = T287 & T286;
  assign T286 = s2_sc_fail ^ 1'h1;
  assign T287 = s2_valid_masked | s2_replay;
  assign T288 = s1_clk_en & T289;
  assign T289 = T304 | T290;
  assign T290 = T299 & T291;
  assign T291 = T296 | T292;
  assign T292 = T295 | T293;
  assign T293 = s4_req_cmd == 5'h4;
  assign T294 = T204 ? s3_req_cmd : s4_req_cmd;
  assign T295 = s4_req_cmd[2'h3];
  assign T296 = T298 | T297;
  assign T297 = s4_req_cmd == 5'h7;
  assign T298 = s4_req_cmd == 5'h1;
  assign T299 = s4_valid & T300;
  assign T300 = T585 == T301;
  assign T301 = s4_req_addr >> 2'h3;
  assign T302 = T204 ? s3_req_addr : s4_req_addr;
  assign T585 = {8'h0, T303};
  assign T303 = s1_addr >> 2'h3;
  assign T586 = reset ? 1'h0 : s3_valid;
  assign T304 = T273 | T259;
  assign T305 = T288 ? 1'h1 : T306;
  assign T306 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T307 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T308 = s2_recycle ? s2_req_typ : T309;
  assign T309 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T310;
  assign T310 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T587 = s2_req_addr[3'h5:1'h0];
  assign T311 = {s3_req_data, s3_req_data};
  assign rowWMask = 1'h1 << rowIdx;
  assign rowIdx = T312;
  assign T312 = s3_req_addr[2'h3];
  assign T588 = s3_req_addr[4'hb:1'h0];
  assign T313 = T249 ? s2_tag_match_way : s3_way;
  assign T314 = T316 & T315;
  assign T315 = FlowThroughSerializer_io_out_bits_client_xact_id < 6'h2;
  assign T316 = FlowThroughSerializer_io_out_valid & T317;
  assign T317 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T321 : T318;
  assign T318 = T320 | T319;
  assign T319 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T320 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T321 = T323 | T322;
  assign T322 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T323 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T324 = T325 | T8;
  assign T325 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T589 = s2_req_addr[4'hb:1'h0];
  assign T590 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T591 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T326 = T327;
  assign T327 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T592 = T328[3'h5:1'h0];
  assign T328 = s2_req_addr >> 3'h6;
  assign T593 = T329[3'h5:1'h0];
  assign T329 = io_cpu_req_bits_addr >> 3'h6;
  assign T330 = s2_recycle ? s2_req_phys : T331;
  assign T331 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T332;
  assign T332 = prober_io_meta_read_valid ? 1'h1 : T333;
  assign T333 = wb_io_meta_read_valid ? 1'h1 : T334;
  assign T334 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T335 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T336 = s1_req_addr >> 4'hc;
  assign T337 = T339 & T338;
  assign T338 = s1_req_phys ^ 1'h1;
  assign T339 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T343 | T340;
  assign T340 = T342 | T341;
  assign T341 = s1_req_cmd == 5'h3;
  assign T342 = s1_req_cmd == 5'h2;
  assign T343 = s1_read | s1_write;
  assign s1_read = T347 | T344;
  assign T344 = T346 | T345;
  assign T345 = s1_req_cmd == 5'h4;
  assign T346 = s1_req_cmd[2'h3];
  assign T347 = T349 | T348;
  assign T348 = s1_req_cmd == 5'h7;
  assign T349 = T351 | T350;
  assign T350 = s1_req_cmd == 5'h6;
  assign T351 = s1_req_cmd == 5'h0;
  assign T352 = T8 & FlowThroughSerializer_io_out_valid;
  assign T353 = cache_pass ^ 1'h1;
  assign cache_pass = T354 | s2_replay;
  assign T354 = s2_valid | s2_killed;
  assign T355 = s1_valid & io_cpu_req_bits_kill;
  assign T356 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R357;
  assign T358 = s1_clk_en ? T359 : R357;
  assign T359 = R360[1'h1:1'h0];
  assign T594 = reset ? 16'h1 : T361;
  assign T361 = T371 ? T362 : R360;
  assign T362 = {T364, T363};
  assign T363 = R360[4'hf:1'h1];
  assign T364 = T366 ^ T365;
  assign T365 = R360[3'h5];
  assign T366 = T368 ^ T367;
  assign T367 = R360[2'h3];
  assign T368 = T370 ^ T369;
  assign T369 = R360[2'h2];
  assign T370 = R360[1'h0];
  assign T371 = T372;
  assign T372 = mshrs_io_req_ready & T431;
  assign T373 = s2_tag_match ? T419 : T374;
  assign T374 = T375[1'h1:1'h0];
  assign T375 = T387 | T376;
  assign T376 = T386 ? T377 : 22'h0;
  assign T377 = T378;
  assign T378 = {R384, R379};
  assign T380 = T381 ? meta_io_resp_3_coh_state : R379;
  assign T381 = s1_clk_en & T382;
  assign T382 = s1_replaced_way_en[2'h3];
  assign s1_replaced_way_en = 1'h1 << T383;
  assign T383 = R360[1'h1:1'h0];
  assign T385 = T381 ? meta_io_resp_3_tag : R384;
  assign T386 = s2_replaced_way_en[2'h3];
  assign T387 = T398 | T388;
  assign T388 = T397 ? T389 : 22'h0;
  assign T389 = T390;
  assign T390 = {R395, R391};
  assign T392 = T393 ? meta_io_resp_2_coh_state : R391;
  assign T393 = s1_clk_en & T394;
  assign T394 = s1_replaced_way_en[2'h2];
  assign T396 = T393 ? meta_io_resp_2_tag : R395;
  assign T397 = s2_replaced_way_en[2'h2];
  assign T398 = T409 | T399;
  assign T399 = T408 ? T400 : 22'h0;
  assign T400 = T401;
  assign T401 = {R406, R402};
  assign T403 = T404 ? meta_io_resp_1_coh_state : R402;
  assign T404 = s1_clk_en & T405;
  assign T405 = s1_replaced_way_en[1'h1];
  assign T407 = T404 ? meta_io_resp_1_tag : R406;
  assign T408 = s2_replaced_way_en[1'h1];
  assign T409 = T418 ? T410 : 22'h0;
  assign T410 = T411;
  assign T411 = {R416, R412};
  assign T413 = T414 ? meta_io_resp_0_coh_state : R412;
  assign T414 = s1_clk_en & T415;
  assign T415 = s1_replaced_way_en[1'h0];
  assign T417 = T414 ? meta_io_resp_0_tag : R416;
  assign T418 = s2_replaced_way_en[1'h0];
  assign T419 = T44;
  assign T420 = s2_tag_match ? T422 : T421;
  assign T421 = T375[5'h15:2'h2];
  assign T422 = T421;
  assign T423 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T424 = s2_recycle ? s2_req_kill : T425;
  assign T425 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T426;
  assign T426 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T427 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T428 = s2_recycle ? s2_req_tag : T429;
  assign T429 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T430;
  assign T430 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T431 = s2_nack_hit ? 1'h0 : T432;
  assign T432 = T454 & T433;
  assign T433 = T441 | T434;
  assign T434 = T438 | T435;
  assign T435 = T437 | T436;
  assign T436 = s2_req_cmd == 5'h4;
  assign T437 = s2_req_cmd[2'h3];
  assign T438 = T440 | T439;
  assign T439 = s2_req_cmd == 5'h7;
  assign T440 = s2_req_cmd == 5'h1;
  assign T441 = T451 | T442;
  assign T442 = T446 | T443;
  assign T443 = T445 | T444;
  assign T444 = s2_req_cmd == 5'h4;
  assign T445 = s2_req_cmd[2'h3];
  assign T446 = T448 | T447;
  assign T447 = s2_req_cmd == 5'h7;
  assign T448 = T450 | T449;
  assign T449 = s2_req_cmd == 5'h6;
  assign T450 = s2_req_cmd == 5'h0;
  assign T451 = T453 | T452;
  assign T452 = s2_req_cmd == 5'h3;
  assign T453 = s2_req_cmd == 5'h2;
  assign T454 = s2_valid_masked & T455;
  assign T455 = s2_hit ^ 1'h1;
  assign T456 = io_mem_probe_valid & T457;
  assign T457 = lrsc_valid ^ 1'h1;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_probe_ready = T458;
  assign T458 = prober_io_req_ready & T459;
  assign T459 = lrsc_valid ^ 1'h1;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_ordered = T460;
  assign T460 = T462 & T461;
  assign T461 = s2_valid ^ 1'h1;
  assign T462 = mshrs_io_fence_rdy & T463;
  assign T463 = s1_valid ^ 1'h1;
  assign io_cpu_xcpt_pf_st = T464;
  assign T464 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T465;
  assign T465 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T466;
  assign T466 = s1_write & misaligned;
  assign misaligned = T467 != 40'h0;
  assign T467 = s1_req_addr & T595;
  assign T595 = {37'h0, T468};
  assign T468 = T469[2'h2:1'h0];
  assign T469 = T470 - 4'h1;
  assign T470 = 1'h1 << T471;
  assign T471 = s1_req_typ[1'h1:1'h0];
  assign io_cpu_xcpt_ma_ld = T472;
  assign T472 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T473;
  assign T473 = s1_replay & s1_read;
  assign io_cpu_resp_bits_store_data = T474;
  assign T474 = cache_pass ? cache_resp_bits_store_data : uncache_resp_bits_store_data;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign cache_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_data_word_bypass = T475;
  assign T475 = {T480, T476};
  assign T476 = T479 ? T478 : T477;
  assign T477 = s2_data_word[5'h1f:1'h0];
  assign T478 = s2_data_word[6'h3f:6'h20];
  assign T479 = s2_req_addr[2'h2];
  assign T480 = T487 ? T482 : T481;
  assign T481 = s2_data_word[6'h3f:6'h20];
  assign T482 = 32'h0 - T596;
  assign T596 = {31'h0, T483};
  assign T483 = T485 & T484;
  assign T484 = T476[5'h1f];
  assign T485 = $signed(1'h0) <= $signed(T486);
  assign T486 = s2_req_typ;
  assign T487 = T488 == 2'h2;
  assign T488 = s2_req_typ[1'h1:1'h0];
  assign io_cpu_resp_bits_has_data = T489;
  assign T489 = cache_pass ? cache_resp_bits_has_data : uncache_resp_bits_has_data;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign cache_resp_bits_has_data = T490;
  assign T490 = T494 | T491;
  assign T491 = T493 | T492;
  assign T492 = s2_req_cmd == 5'h4;
  assign T493 = s2_req_cmd[2'h3];
  assign T494 = T496 | T495;
  assign T495 = s2_req_cmd == 5'h7;
  assign T496 = T498 | T497;
  assign T497 = s2_req_cmd == 5'h6;
  assign T498 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_replay = T499;
  assign T499 = cache_pass ? cache_resp_bits_replay : uncache_resp_bits_replay;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign cache_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T500;
  assign T500 = cache_pass ? cache_resp_bits_nack : uncache_resp_bits_nack;
  assign uncache_resp_bits_nack = mshrs_io_resp_bits_nack;
  assign cache_resp_bits_nack = T501;
  assign T501 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T502;
  assign T502 = cache_pass ? cache_resp_bits_data : uncache_resp_bits_data;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign cache_resp_bits_data = T503;
  assign T503 = T504 | T597;
  assign T597 = {63'h0, s2_sc_fail};
  assign T504 = {T532, T505};
  assign T505 = s2_sc ? 8'h0 : T506;
  assign T506 = T531 ? T530 : T507;
  assign T507 = T508[3'h7:1'h0];
  assign T508 = {T524, T509};
  assign T509 = T523 ? T522 : T510;
  assign T510 = T511[4'hf:1'h0];
  assign T511 = {T516, T512};
  assign T512 = T515 ? T514 : T513;
  assign T513 = s2_data_word[5'h1f:1'h0];
  assign T514 = s2_data_word[6'h3f:6'h20];
  assign T515 = s2_req_addr[2'h2];
  assign T516 = T521 ? T518 : T517;
  assign T517 = s2_data_word[6'h3f:6'h20];
  assign T518 = 32'h0 - T598;
  assign T598 = {31'h0, T519};
  assign T519 = T485 & T520;
  assign T520 = T512[5'h1f];
  assign T521 = T488 == 2'h2;
  assign T522 = T511[5'h1f:5'h10];
  assign T523 = s2_req_addr[1'h1];
  assign T524 = T529 ? T526 : T525;
  assign T525 = T511[6'h3f:5'h10];
  assign T526 = 48'h0 - T599;
  assign T599 = {47'h0, T527};
  assign T527 = T485 & T528;
  assign T528 = T509[4'hf];
  assign T529 = T488 == 2'h1;
  assign T530 = T508[4'hf:4'h8];
  assign T531 = s2_req_addr[1'h0];
  assign T532 = T537 ? T534 : T533;
  assign T533 = T508[6'h3f:4'h8];
  assign T534 = 56'h0 - T600;
  assign T600 = {55'h0, T535};
  assign T535 = T485 & T536;
  assign T536 = T505[3'h7];
  assign T537 = T538 | s2_sc;
  assign T538 = T488 == 2'h0;
  assign io_cpu_resp_bits_typ = T539;
  assign T539 = cache_pass ? cache_resp_bits_typ : uncache_resp_bits_typ;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign cache_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_cmd = T540;
  assign T540 = cache_pass ? cache_resp_bits_cmd : uncache_resp_bits_cmd;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_tag = T541;
  assign T541 = cache_pass ? cache_resp_bits_tag : uncache_resp_bits_tag;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign cache_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_addr = T542;
  assign T542 = cache_pass ? cache_resp_bits_addr : uncache_resp_bits_addr;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign cache_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_valid = T543;
  assign T543 = cache_pass ? cache_resp_valid : uncache_resp_valid;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign cache_resp_valid = T544;
  assign T544 = T546 & T545;
  assign T545 = s2_data_correctable ^ 1'h1;
  assign T546 = s2_replay | T547;
  assign T547 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T548;
  assign T548 = block_miss ? 1'h0 : T549;
  assign T549 = T556 ? 1'h0 : T550;
  assign T550 = T555 ? 1'h0 : T551;
  assign T551 = T552 == 1'h0;
  assign T552 = T554 & T553;
  assign T553 = io_cpu_req_bits_phys ^ 1'h1;
  assign T554 = dtlb_io_req_ready ^ 1'h1;
  assign T555 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T556 = readArb_io_in_3_ready ^ 1'h1;
  assign T601 = reset ? 1'h0 : T557;
  assign T557 = T558 & s2_nack_miss;
  assign T558 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_req_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_req_bits_data( wbArb_io_out_bits_data ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       //.io_meta_read_bits_way_en(  )
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_release_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_release_bits_r_type( wb_io_release_bits_r_type ),
       .io_release_bits_data( wb_io_release_bits_data )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T456 ),
       .io_req_bits_addr_block( io_mem_probe_bits_addr_block ),
       .io_req_bits_p_type( io_mem_probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_rep_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       //.io_meta_read_bits_way_en(  )
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( prober_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_block_state_state( T44 )
  );
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T431 ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T420 ),
       .io_req_bits_old_meta_coh_state( T373 ),
       .io_req_bits_way_en( T356 ),
       .io_resp_ready( T353 ),
       .io_resp_valid( mshrs_io_resp_valid ),
       .io_resp_bits_addr( mshrs_io_resp_bits_addr ),
       .io_resp_bits_tag( mshrs_io_resp_bits_tag ),
       .io_resp_bits_cmd( mshrs_io_resp_bits_cmd ),
       .io_resp_bits_typ( mshrs_io_resp_bits_typ ),
       .io_resp_bits_data( mshrs_io_resp_bits_data ),
       .io_resp_bits_nack( mshrs_io_resp_bits_nack ),
       .io_resp_bits_replay( mshrs_io_resp_bits_replay ),
       .io_resp_bits_has_data( mshrs_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( mshrs_io_resp_bits_store_data ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( io_mem_acquire_ready ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( mshrs_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( mshrs_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( mshrs_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( mshrs_io_mem_req_bits_union ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_refill_way_en( mshrs_io_refill_way_en ),
       .io_refill_addr( mshrs_io_refill_addr ),
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       .io_meta_read_bits_way_en( mshrs_io_meta_read_bits_way_en ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T352 ),
       .io_mem_grant_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_mem_grant_bits_data( FlowThroughSerializer_io_out_bits_data ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( mshrs_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T337 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T336 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_req_bits_store( s1_write ),
       .io_resp_miss( dtlb_io_resp_miss ),
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dtlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dtlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dtlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dtlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_read_bits_way_en( metaReadArb_io_out_bits_way_en ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_3_tag( meta_io_resp_3_tag ),
       .io_resp_3_coh_state( meta_io_resp_3_coh_state ),
       .io_resp_2_tag( meta_io_resp_2_tag ),
       .io_resp_2_coh_state( meta_io_resp_2_coh_state ),
       .io_resp_1_tag( meta_io_resp_1_tag ),
       .io_resp_1_coh_state( meta_io_resp_1_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state ),
       .init( init )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T593 ),
       //.io_in_4_bits_way_en(  )
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       //.io_in_3_bits_way_en(  )
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       //.io_in_2_bits_way_en(  )
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_meta_read_bits_way_en ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T592 ),
       //.io_in_0_bits_way_en(  )
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaReadArb_io_out_bits_way_en )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign metaReadArb.io_in_4_bits_way_en = {1{$random}};
    assign metaReadArb.io_in_3_bits_way_en = {1{$random}};
    assign metaReadArb.io_in_2_bits_way_en = {1{$random}};
    assign metaReadArb.io_in_0_bits_way_en = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T326 ),
       .io_resp_3( data_io_resp_3 ),
       .io_resp_2( data_io_resp_2 ),
       .io_resp_1( data_io_resp_1 ),
       .io_resp_0( data_io_resp_0 ),
       .init( init )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 4'hf ),
       .io_in_3_bits_addr( T591 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 4'hf ),
       .io_in_1_bits_addr( T590 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 4'hf ),
       .io_in_0_bits_addr( T589 ),
       .io_out_ready( T324 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T314 ),
       .io_in_1_bits_way_en( mshrs_io_refill_way_en ),
       .io_in_1_bits_addr( mshrs_io_refill_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( FlowThroughSerializer_io_out_bits_data ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T588 ),
       .io_in_0_bits_wmask( rowWMask ),
       .io_in_0_bits_data( T311 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T587 ),
       .io_cmd( s2_req_cmd ),
       .io_typ( s2_req_typ ),
       .io_lhs( T568 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  LockingArbiter_0 releaseArb(.clk(clk), .reset(reset),
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_in_1_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_in_0_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_out_ready( io_mem_release_ready ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr_beat( releaseArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( releaseArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( releaseArb_io_out_bits_voluntary ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type ),
       .io_out_bits_data( releaseArb_io_out_bits_data )
       //.io_chosen(  )
  );
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( T8 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_1_bits_data( mshrs_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_in_0_bits_data( prober_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_out_bits_data( wbArb_io_out_bits_data ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "DCache exception occurred - cache response not killed.");
    $finish;
  end
// synthesis translate_on
`endif
    R4 <= T5;
    if(T138) begin
      s2_req_data <= s1_req_data;
    end else if(T21) begin
      s2_req_data <= T19;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T20;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T30) begin
      s2_recycle_next <= s2_recycle_ecc;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T31;
    end
    if(s1_clk_en) begin
      R48 <= meta_io_resp_3_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T563;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T562;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T564;
    end
    if(s1_clk_en) begin
      R92 <= meta_io_resp_2_coh_state;
    end
    if(s1_clk_en) begin
      R98 <= meta_io_resp_1_coh_state;
    end
    if(s1_clk_en) begin
      R103 <= meta_io_resp_0_coh_state;
    end
    if(reset) begin
      R129 <= 1'h0;
    end else begin
      R129 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R145 <= T569;
    if(T153) begin
      R150 <= T152;
    end
    R162 <= T571;
    if(T170) begin
      R167 <= T169;
    end
    R176 <= T573;
    if(T184) begin
      R181 <= T183;
    end
    R189 <= T575;
    if(T197) begin
      R194 <= T196;
    end
    if(T288) begin
      s2_store_bypass_data <= T201;
    end
    if(T204) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T205;
    end
    if(T220) begin
      lrsc_addr <= T219;
    end
    if(T234) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_invalidate_lr) begin
      lrsc_count <= 5'h0;
    end else if(T242) begin
      lrsc_count <= 5'h0;
    end else if(T240) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T239;
    end
    s3_req_data <= T580;
    if(T249) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T249) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T204) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T204) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T288) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T249) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    s2_killed <= T355;
    if(s1_clk_en) begin
      R357 <= T359;
    end
    if(reset) begin
      R360 <= 16'h1;
    end else if(T371) begin
      R360 <= T362;
    end
    if(T381) begin
      R379 <= meta_io_resp_3_coh_state;
    end
    if(T381) begin
      R384 <= meta_io_resp_3_tag;
    end
    if(T393) begin
      R391 <= meta_io_resp_2_coh_state;
    end
    if(T393) begin
      R395 <= meta_io_resp_2_tag;
    end
    if(T404) begin
      R402 <= meta_io_resp_1_coh_state;
    end
    if(T404) begin
      R406 <= meta_io_resp_1_tag;
    end
    if(T414) begin
      R412 <= meta_io_resp_0_coh_state;
    end
    if(T414) begin
      R416 <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T557;
    end
  end
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [26:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_prv,
    input  io_in_1_bits_store,
    input  io_in_1_bits_fetch,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [26:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_prv,
    input  io_in_0_bits_store,
    input  io_in_0_bits_fetch,
    input  io_out_ready,
    output io_out_valid,
    output[26:0] io_out_bits_addr,
    output[1:0] io_out_bits_prv,
    output io_out_bits_store,
    output io_out_bits_fetch,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T28;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire[26:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T28 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_fetch = T5;
  assign T5 = T6 ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T6 = chosen;
  assign io_out_bits_store = T7;
  assign T7 = T6 ? io_in_1_bits_store : io_in_0_bits_store;
  assign io_out_bits_prv = T8;
  assign T8 = T6 ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign io_out_bits_addr = T9;
  assign T9 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = last_grant < 1'h0;
  assign T19 = last_grant < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = last_grant < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [26:0] io_requestor_1_req_bits_addr,
    input [1:0] io_requestor_1_req_bits_prv,
    input  io_requestor_1_req_bits_store,
    input  io_requestor_1_req_bits_fetch,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[19:0] io_requestor_1_resp_bits_pte_ppn,
    output[2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
    output io_requestor_1_resp_bits_pte_d,
    output io_requestor_1_resp_bits_pte_r,
    output[3:0] io_requestor_1_resp_bits_pte_typ,
    output io_requestor_1_resp_bits_pte_v,
    output io_requestor_1_status_sd,
    output[30:0] io_requestor_1_status_zero2,
    output io_requestor_1_status_sd_rv32,
    output[8:0] io_requestor_1_status_zero1,
    output[4:0] io_requestor_1_status_vm,
    output io_requestor_1_status_mprv,
    output[1:0] io_requestor_1_status_xs,
    output[1:0] io_requestor_1_status_fs,
    output[1:0] io_requestor_1_status_prv3,
    output io_requestor_1_status_ie3,
    output[1:0] io_requestor_1_status_prv2,
    output io_requestor_1_status_ie2,
    output[1:0] io_requestor_1_status_prv1,
    output io_requestor_1_status_ie1,
    output[1:0] io_requestor_1_status_prv,
    output io_requestor_1_status_ie,
    output io_requestor_1_invalidate,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [26:0] io_requestor_0_req_bits_addr,
    input [1:0] io_requestor_0_req_bits_prv,
    input  io_requestor_0_req_bits_store,
    input  io_requestor_0_req_bits_fetch,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[19:0] io_requestor_0_resp_bits_pte_ppn,
    output[2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
    output io_requestor_0_resp_bits_pte_d,
    output io_requestor_0_resp_bits_pte_r,
    output[3:0] io_requestor_0_resp_bits_pte_typ,
    output io_requestor_0_resp_bits_pte_v,
    output io_requestor_0_status_sd,
    output[30:0] io_requestor_0_status_zero2,
    output io_requestor_0_status_sd_rv32,
    output[8:0] io_requestor_0_status_zero1,
    output[4:0] io_requestor_0_status_vm,
    output io_requestor_0_status_mprv,
    output[1:0] io_requestor_0_status_xs,
    output[1:0] io_requestor_0_status_fs,
    output[1:0] io_requestor_0_status_prv3,
    output io_requestor_0_status_ie3,
    output[1:0] io_requestor_0_status_prv2,
    output io_requestor_0_status_ie2,
    output[1:0] io_requestor_0_status_prv1,
    output io_requestor_0_status_ie1,
    output[1:0] io_requestor_0_status_prv,
    output io_requestor_0_status_ie,
    output io_requestor_0_invalidate,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    //output[9:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [9:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [9:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_status_sd,
    input [30:0] io_dpath_status_zero2,
    input  io_dpath_status_sd_rv32,
    input [8:0] io_dpath_status_zero1,
    input [4:0] io_dpath_status_vm,
    input  io_dpath_status_mprv,
    input [1:0] io_dpath_status_xs,
    input [1:0] io_dpath_status_fs,
    input [1:0] io_dpath_status_prv3,
    input  io_dpath_status_ie3,
    input [1:0] io_dpath_status_prv2,
    input  io_dpath_status_ie2,
    input [1:0] io_dpath_status_prv1,
    input  io_dpath_status_ie1,
    input [1:0] io_dpath_status_prv,
    input  io_dpath_status_ie
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T227;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] count;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire pte_cache_hit;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[1:0] T26;
  reg  R27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T228;
  wire[1:0] T229;
  wire T230;
  wire[2:0] T36;
  wire T231;
  wire[1:0] T37;
  wire[2:0] T38;
  wire T39;
  reg [2:0] R40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire[2:0] T44;
  wire[5:0] T45;
  wire[1:0] T46;
  wire T47;
  wire[1:0] T232;
  wire T233;
  wire[1:0] T234;
  wire[1:0] T235;
  wire T236;
  wire T237;
  wire T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  reg  R68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire T81;
  wire[31:0] pte_addr;
  wire[28:0] T82;
  wire[28:0] T83;
  wire[8:0] vpn_idx;
  wire[8:0] T84;
  wire[8:0] T85;
  wire[8:0] T86;
  reg [26:0] r_req_addr;
  wire[26:0] T87;
  wire T88;
  wire[8:0] T89;
  wire[17:0] T90;
  wire T91;
  wire[1:0] T92;
  wire[8:0] T93;
  wire[26:0] T94;
  wire T95;
  reg [19:0] r_pte_ppn;
  wire[19:0] T96;
  wire[19:0] T97;
  wire[19:0] T98;
  wire[19:0] T99;
  wire[19:0] T100;
  wire T101;
  wire T102;
  wire set_dirty_bit;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  reg  r_req_store;
  wire T107;
  wire T108;
  wire T109;
  wire perm_ok;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  reg  r_req_fetch;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  reg [1:0] r_req_prv;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire[19:0] pte_cache_data;
  wire[19:0] T145;
  wire[19:0] T146;
  reg [19:0] T147 [2:0];
  wire[19:0] T148;
  wire T149;
  wire T150;
  wire[1:0] T151;
  wire T152;
  wire[19:0] T153;
  wire[19:0] T154;
  wire[19:0] T155;
  wire T156;
  wire[19:0] T157;
  wire[19:0] T158;
  wire T159;
  wire[31:0] T160;
  reg [31:0] T161 [2:0];
  wire[31:0] T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire[31:0] T167;
  wire T168;
  wire[31:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[2:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire[63:0] T238;
  wire[29:0] T193;
  wire[29:0] T194;
  wire[5:0] T195;
  wire[4:0] T196;
  wire pte_wdata_v;
  wire[3:0] pte_wdata_typ;
  wire pte_wdata_r;
  wire[23:0] T197;
  wire[3:0] T198;
  wire pte_wdata_d;
  wire[2:0] pte_wdata_reserved_for_software;
  wire[19:0] pte_wdata_ppn;
  wire[4:0] T199;
  wire T200;
  wire[39:0] T239;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  reg  r_pte_v;
  wire T205;
  reg [3:0] r_pte_typ;
  wire[3:0] T206;
  reg  r_pte_r;
  wire T207;
  reg  r_pte_d;
  wire T208;
  reg [2:0] r_pte_reserved_for_software;
  wire[2:0] T209;
  wire[2:0] T210;
  wire[19:0] T240;
  wire[27:0] resp_ppn;
  wire[27:0] T211;
  wire[27:0] T212;
  wire[17:0] T213;
  wire[9:0] T214;
  wire[27:0] T215;
  wire[8:0] T216;
  wire[18:0] T217;
  wire T218;
  wire[1:0] T219;
  wire[27:0] r_resp_ppn;
  wire T220;
  wire resp_err;
  wire T221;
  wire T222;
  reg  r_req_dest;
  wire T223;
  wire resp_val;
  wire T224;
  wire[19:0] T241;
  wire T225;
  wire T226;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[26:0] arb_io_out_bits_addr;
  wire[1:0] arb_io_out_bits_prv;
  wire arb_io_out_bits_store;
  wire arb_io_out_bits_fetch;
  wire arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    R27 = {1{$random}};
    R40 = {1{$random}};
    R68 = {1{$random}};
    R73 = {1{$random}};
    r_req_addr = {1{$random}};
    r_pte_ppn = {1{$random}};
    r_req_store = {1{$random}};
    r_req_fetch = {1{$random}};
    r_req_prv = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T147[initvar] = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T161[initvar] = {1{$random}};
    r_pte_v = {1{$random}};
    r_pte_typ = {1{$random}};
    r_pte_r = {1{$random}};
    r_pte_d = {1{$random}};
    r_pte_reserved_for_software = {1{$random}};
    r_req_dest = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
//  assign io_mem_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = state == 3'h0;
  assign T227 = reset ? 3'h0 : T1;
  assign T1 = T192 ? 3'h0 : T2;
  assign T2 = T191 ? 3'h0 : T3;
  assign T3 = T190 ? 3'h1 : T4;
  assign T4 = T188 ? 3'h3 : T5;
  assign T5 = T186 ? 3'h4 : T6;
  assign T6 = T183 ? T182 : T7;
  assign T7 = T177 ? 3'h1 : T8;
  assign T8 = T176 ? 3'h6 : T9;
  assign T9 = T174 ? 3'h1 : T10;
  assign T10 = T171 ? 3'h2 : T11;
  assign T11 = T15 ? 3'h1 : T12;
  assign T12 = T13 ? 3'h1 : state;
  assign T13 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T15 = T170 & T16;
  assign T16 = pte_cache_hit & T17;
  assign T17 = count < 2'h2;
  assign T18 = T177 ? T22 : T19;
  assign T19 = T15 ? T21 : T20;
  assign T20 = T14 ? 2'h0 : count;
  assign T21 = count + 2'h1;
  assign T22 = count + 2'h1;
  assign pte_cache_hit = T23 != 3'h0;
  assign T23 = T78 & T24;
  assign T24 = T25;
  assign T25 = {R73, T26};
  assign T26 = {R68, R27};
  assign T28 = T67 ? 1'h0 : T29;
  assign T29 = T30 ? 1'h1 : R27;
  assign T30 = T60 & T31;
  assign T31 = T32[1'h0];
  assign T32 = 1'h1 << T33;
  assign T33 = T34;
  assign T34 = T59 ? T37 : T228;
  assign T228 = T231 ? 1'h0 : T229;
  assign T229 = T230 ? 1'h1 : 2'h2;
  assign T230 = T36[1'h1];
  assign T36 = ~ T24;
  assign T231 = T36[1'h0];
  assign T37 = T38[1'h1:1'h0];
  assign T38 = {T57, T39};
  assign T39 = R40[T57];
  assign T41 = T55 ? T42 : R40;
  assign T42 = T50 | T43;
  assign T43 = T49 ? 3'h0 : T44;
  assign T44 = T45[2'h2:1'h0];
  assign T45 = 3'h1 << T46;
  assign T46 = {1'h1, T47};
  assign T47 = T232[1'h1];
  assign T232 = {T237, T233};
  assign T233 = T234[1'h1];
  assign T234 = T236 | T235;
  assign T235 = T23[1'h1:1'h0];
  assign T236 = T23[2'h2];
  assign T237 = T236 != 1'h0;
  assign T49 = T232[1'h0];
  assign T50 = T52 & T51;
  assign T51 = ~ T44;
  assign T52 = T54 | T53;
  assign T53 = T47 ? 3'h0 : 3'h2;
  assign T54 = R40 & 3'h5;
  assign T55 = pte_cache_hit & T56;
  assign T56 = state == 3'h1;
  assign T57 = {1'h1, T58};
  assign T58 = R40[1'h1];
  assign T59 = T24 == 3'h7;
  assign T60 = T62 & T61;
  assign T61 = pte_cache_hit ^ 1'h1;
  assign T62 = io_mem_resp_valid & T63;
  assign T63 = T66 & T64;
  assign T64 = T65 < 4'h2;
  assign T65 = io_mem_resp_bits_data[3'h4:1'h1];
  assign T66 = io_mem_resp_bits_data[1'h0];
  assign T67 = reset | io_dpath_invalidate;
  assign T69 = T67 ? 1'h0 : T70;
  assign T70 = T71 ? 1'h1 : R68;
  assign T71 = T60 & T72;
  assign T72 = T32[1'h1];
  assign T74 = T67 ? 1'h0 : T75;
  assign T75 = T76 ? 1'h1 : R73;
  assign T76 = T60 & T77;
  assign T77 = T32[2'h2];
  assign T78 = T79;
  assign T79 = {T168, T80};
  assign T80 = {T166, T81};
  assign T81 = T160 == pte_addr;
  assign pte_addr = T82 << 2'h3;
  assign T82 = T83;
  assign T83 = {r_pte_ppn, vpn_idx};
  assign vpn_idx = T95 ? T93 : T84;
  assign T84 = T91 ? T89 : T85;
  assign T85 = T86;
  assign T86 = r_req_addr >> 5'h12;
  assign T87 = T88 ? arb_io_out_bits_addr : r_req_addr;
  assign T88 = T0 & arb_io_out_valid;
  assign T89 = T90[4'h8:1'h0];
  assign T90 = r_req_addr >> 4'h9;
  assign T91 = T92[1'h0];
  assign T92 = count;
  assign T93 = T94[4'h8:1'h0];
  assign T94 = r_req_addr >> 1'h0;
  assign T95 = T92[1'h1];
  assign T96 = T15 ? pte_cache_data : T97;
  assign T97 = T101 ? T100 : T98;
  assign T98 = T88 ? T99 : r_pte_ppn;
  assign T99 = io_dpath_ptbr[5'h1f:4'hc];
  assign T100 = io_mem_resp_bits_data[5'h1d:4'ha];
  assign T101 = T143 & T102;
  assign T102 = set_dirty_bit ^ 1'h1;
  assign set_dirty_bit = perm_ok & T103;
  assign T103 = T108 | T104;
  assign T104 = r_req_store & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = io_mem_resp_bits_data[3'h6];
  assign T107 = T88 ? arb_io_out_bits_store : r_req_store;
  assign T108 = T109 ^ 1'h1;
  assign T109 = io_mem_resp_bits_data[3'h5];
  assign perm_ok = T141 ? T129 : T110;
  assign T110 = r_req_fetch ? T122 : T111;
  assign T111 = r_req_store ? T116 : T112;
  assign T112 = T114 & T113;
  assign T113 = T65 < 4'h8;
  assign T114 = T66 & T115;
  assign T115 = 4'h2 <= T65;
  assign T116 = T118 & T117;
  assign T117 = T65[1'h0];
  assign T118 = T120 & T119;
  assign T119 = T65 < 4'h8;
  assign T120 = T66 & T121;
  assign T121 = 4'h2 <= T65;
  assign T122 = T124 & T123;
  assign T123 = T65[1'h1];
  assign T124 = T126 & T125;
  assign T125 = T65 < 4'h8;
  assign T126 = T66 & T127;
  assign T127 = 4'h2 <= T65;
  assign T128 = T88 ? arb_io_out_bits_fetch : r_req_fetch;
  assign T129 = r_req_fetch ? T137 : T130;
  assign T130 = r_req_store ? T133 : T131;
  assign T131 = T66 & T132;
  assign T132 = 4'h2 <= T65;
  assign T133 = T135 & T134;
  assign T134 = T65[1'h0];
  assign T135 = T66 & T136;
  assign T136 = 4'h2 <= T65;
  assign T137 = T139 & T138;
  assign T138 = T65[1'h1];
  assign T139 = T66 & T140;
  assign T140 = 4'h4 <= T65;
  assign T141 = r_req_prv[1'h0];
  assign T142 = T88 ? arb_io_out_bits_prv : r_req_prv;
  assign T143 = io_mem_resp_valid & T144;
  assign T144 = state == 3'h2;
  assign pte_cache_data = T153 | T145;
  assign T145 = T152 ? T146 : 20'h0;
  assign T146 = T147[2'h2];
  assign T149 = T60 & T150;
  assign T150 = T151 < 2'h3;
  assign T151 = T34;
  assign T152 = T23[2'h2];
  assign T153 = T157 | T154;
  assign T154 = T156 ? T155 : 20'h0;
  assign T155 = T147[2'h1];
  assign T156 = T23[1'h1];
  assign T157 = T159 ? T158 : 20'h0;
  assign T158 = T147[2'h0];
  assign T159 = T23[1'h0];
  assign T160 = T161[2'h0];
  assign T163 = T60 & T164;
  assign T164 = T165 < 2'h3;
  assign T165 = T34;
  assign T166 = T167 == pte_addr;
  assign T167 = T161[2'h1];
  assign T168 = T169 == pte_addr;
  assign T169 = T161[2'h2];
  assign T170 = 3'h1 == state;
  assign T171 = T170 & T172;
  assign T172 = T173 & io_mem_req_ready;
  assign T173 = T16 ^ 1'h1;
  assign T174 = T175 & io_mem_resp_bits_nack;
  assign T175 = 3'h2 == state;
  assign T176 = T175 & io_mem_resp_valid;
  assign T177 = T176 & T178;
  assign T178 = T180 & T179;
  assign T179 = count < 2'h2;
  assign T180 = T66 & T181;
  assign T181 = T65 < 4'h2;
  assign T182 = set_dirty_bit ? 3'h3 : 3'h5;
  assign T183 = T176 & T184;
  assign T184 = T66 & T185;
  assign T185 = 4'h2 <= T65;
  assign T186 = T187 & io_mem_req_ready;
  assign T187 = 3'h3 == state;
  assign T188 = T189 & io_mem_resp_bits_nack;
  assign T189 = 3'h4 == state;
  assign T190 = T189 & io_mem_resp_valid;
  assign T191 = 3'h5 == state;
  assign T192 = 3'h6 == state;
  assign io_mem_req_bits_data = T238;
  assign T238 = {34'h0, T193};
  assign T193 = T194;
  assign T194 = {T197, T195};
  assign T195 = {pte_wdata_r, T196};
  assign T196 = {pte_wdata_typ, pte_wdata_v};
  assign pte_wdata_v = 1'h0;
  assign pte_wdata_typ = 4'h0;
  assign pte_wdata_r = 1'h1;
  assign T197 = {pte_wdata_ppn, T198};
  assign T198 = {pte_wdata_reserved_for_software, pte_wdata_d};
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_reserved_for_software = 3'h0;
  assign pte_wdata_ppn = 20'h0;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_cmd = T199;
  assign T199 = T200 ? 5'ha : 5'h0;
  assign T200 = state == 3'h3;
  assign io_mem_req_bits_addr = T239;
  assign T239 = {8'h0, pte_addr};
  assign io_mem_req_valid = T201;
  assign T201 = T15 ? 1'h0 : T202;
  assign T202 = T204 | T203;
  assign T203 = state == 3'h3;
  assign T204 = state == 3'h1;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_ie = io_dpath_status_ie;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_0_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_0_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_0_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_0_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_0_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign T205 = T101 ? T66 : r_pte_v;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign T206 = T101 ? T65 : r_pte_typ;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign T207 = T101 ? T109 : r_pte_r;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign T208 = T101 ? T106 : r_pte_d;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign T209 = T101 ? T210 : r_pte_reserved_for_software;
  assign T210 = io_mem_resp_bits_data[4'h9:3'h7];
  assign io_requestor_0_resp_bits_pte_ppn = T240;
  assign T240 = resp_ppn[5'h13:1'h0];
  assign resp_ppn = T220 ? r_resp_ppn : T211;
  assign T211 = T218 ? T215 : T212;
  assign T212 = {T214, T213};
  assign T213 = r_req_addr[5'h11:1'h0];
  assign T214 = r_resp_ppn >> 5'h12;
  assign T215 = {T217, T216};
  assign T216 = r_req_addr[4'h8:1'h0];
  assign T217 = r_resp_ppn >> 4'h9;
  assign T218 = T219[1'h0];
  assign T219 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hc;
  assign T220 = T219[1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = state == 3'h6;
  assign io_requestor_0_resp_valid = T221;
  assign T221 = resp_val & T222;
  assign T222 = r_req_dest == 1'h0;
  assign T223 = T88 ? arb_io_chosen : r_req_dest;
  assign resp_val = T224 | resp_err;
  assign T224 = state == 3'h5;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_ie = io_dpath_status_ie;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_1_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_1_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_1_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_1_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_1_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_ppn = T241;
  assign T241 = resp_ppn[5'h13:1'h0];
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T225;
  assign T225 = resp_val & T226;
  assign T226 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_3 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits_addr( io_requestor_1_req_bits_addr ),
       .io_in_1_bits_prv( io_requestor_1_req_bits_prv ),
       .io_in_1_bits_store( io_requestor_1_req_bits_store ),
       .io_in_1_bits_fetch( io_requestor_1_req_bits_fetch ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits_addr( io_requestor_0_req_bits_addr ),
       .io_in_0_bits_prv( io_requestor_0_req_bits_prv ),
       .io_in_0_bits_store( io_requestor_0_req_bits_store ),
       .io_in_0_bits_fetch( io_requestor_0_req_bits_fetch ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits_addr( arb_io_out_bits_addr ),
       .io_out_bits_prv( arb_io_out_bits_prv ),
       .io_out_bits_store( arb_io_out_bits_store ),
       .io_out_bits_fetch( arb_io_out_bits_fetch ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T192) begin
      state <= 3'h0;
    end else if(T191) begin
      state <= 3'h0;
    end else if(T190) begin
      state <= 3'h1;
    end else if(T188) begin
      state <= 3'h3;
    end else if(T186) begin
      state <= 3'h4;
    end else if(T183) begin
      state <= T182;
    end else if(T177) begin
      state <= 3'h1;
    end else if(T176) begin
      state <= 3'h6;
    end else if(T174) begin
      state <= 3'h1;
    end else if(T171) begin
      state <= 3'h2;
    end else if(T15) begin
      state <= 3'h1;
    end else if(T13) begin
      state <= 3'h1;
    end
    if(T177) begin
      count <= T22;
    end else if(T15) begin
      count <= T21;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T67) begin
      R27 <= 1'h0;
    end else if(T30) begin
      R27 <= 1'h1;
    end
    if(T55) begin
      R40 <= T42;
    end
    if(T67) begin
      R68 <= 1'h0;
    end else if(T71) begin
      R68 <= 1'h1;
    end
    if(T67) begin
      R73 <= 1'h0;
    end else if(T76) begin
      R73 <= 1'h1;
    end
    if(T88) begin
      r_req_addr <= arb_io_out_bits_addr;
    end
    if(T15) begin
      r_pte_ppn <= pte_cache_data;
    end else if(T101) begin
      r_pte_ppn <= T100;
    end else if(T88) begin
      r_pte_ppn <= T99;
    end
    if(T88) begin
      r_req_store <= arb_io_out_bits_store;
    end
    if(T88) begin
      r_req_fetch <= arb_io_out_bits_fetch;
    end
    if(T88) begin
      r_req_prv <= arb_io_out_bits_prv;
    end
    if (T149)
      T147[T34] <= T100;
    if (T163)
      T161[T34] <= pte_addr;
    if(T101) begin
      r_pte_v <= T66;
    end
    if(T101) begin
      r_pte_typ <= T65;
    end
    if(T101) begin
      r_pte_r <= T109;
    end
    if(T101) begin
      r_pte_d <= T106;
    end
    if(T101) begin
      r_pte_reserved_for_software <= T210;
    end
    if(T88) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_2_req_ready,
    input  io_requestor_2_req_valid,
    input [39:0] io_requestor_2_req_bits_addr,
    input [9:0] io_requestor_2_req_bits_tag,
    input [4:0] io_requestor_2_req_bits_cmd,
    input [2:0] io_requestor_2_req_bits_typ,
    input  io_requestor_2_req_bits_kill,
    input  io_requestor_2_req_bits_phys,
    input [63:0] io_requestor_2_req_bits_data,
    output io_requestor_2_resp_valid,
    output[39:0] io_requestor_2_resp_bits_addr,
    output[9:0] io_requestor_2_resp_bits_tag,
    output[4:0] io_requestor_2_resp_bits_cmd,
    output[2:0] io_requestor_2_resp_bits_typ,
    output[63:0] io_requestor_2_resp_bits_data,
    output io_requestor_2_resp_bits_nack,
    output io_requestor_2_resp_bits_replay,
    output io_requestor_2_resp_bits_has_data,
    output[63:0] io_requestor_2_resp_bits_data_word_bypass,
    output[63:0] io_requestor_2_resp_bits_store_data,
    output io_requestor_2_replay_next_valid,
    output[9:0] io_requestor_2_replay_next_bits,
    output io_requestor_2_xcpt_ma_ld,
    output io_requestor_2_xcpt_ma_st,
    output io_requestor_2_xcpt_pf_ld,
    output io_requestor_2_xcpt_pf_st,
    //input  io_requestor_2_invalidate_lr
    output io_requestor_2_ordered,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [39:0] io_requestor_1_req_bits_addr,
    input [9:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_kill,
    input  io_requestor_1_req_bits_phys,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[39:0] io_requestor_1_resp_bits_addr,
    output[9:0] io_requestor_1_resp_bits_tag,
    output[4:0] io_requestor_1_resp_bits_cmd,
    output[2:0] io_requestor_1_resp_bits_typ,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_word_bypass,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[9:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    input  io_requestor_1_invalidate_lr,
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [39:0] io_requestor_0_req_bits_addr,
    input [9:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_kill,
    input  io_requestor_0_req_bits_phys,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[39:0] io_requestor_0_resp_bits_addr,
    output[9:0] io_requestor_0_resp_bits_tag,
    output[4:0] io_requestor_0_resp_bits_cmd,
    output[2:0] io_requestor_0_resp_bits_typ,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_word_bypass,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[9:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_invalidate_lr
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    output[9:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [9:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [9:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered
);

  wire[63:0] T0;
  wire[63:0] T1;
  reg  r_valid_1;
  reg  r_valid_0;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[4:0] T8;
  wire[4:0] T9;
  wire[9:0] T53;
  wire[11:0] T10;
  wire[11:0] T11;
  wire[11:0] T12;
  wire[11:0] T13;
  wire[11:0] T14;
  wire[39:0] T15;
  wire[39:0] T16;
  wire T17;
  wire T18;
  wire[9:0] T54;
  wire[7:0] T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire[9:0] T55;
  wire[7:0] T27;
  wire T28;
  wire[9:0] T56;
  wire[7:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire T36;
  wire[9:0] T57;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[9:0] T58;
  wire[7:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire[9:0] T59;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_valid_1 = {1{$random}};
    r_valid_0 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : T1;
  assign T1 = r_valid_1 ? io_requestor_1_req_bits_data : io_requestor_2_req_bits_data;
  assign io_mem_req_bits_phys = T2;
  assign T2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : T3;
  assign T3 = io_requestor_1_req_valid ? io_requestor_1_req_bits_phys : io_requestor_2_req_bits_phys;
  assign io_mem_req_bits_kill = T4;
  assign T4 = r_valid_0 ? io_requestor_0_req_bits_kill : T5;
  assign T5 = r_valid_1 ? io_requestor_1_req_bits_kill : io_requestor_2_req_bits_kill;
  assign io_mem_req_bits_typ = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : T7;
  assign T7 = io_requestor_1_req_valid ? io_requestor_1_req_bits_typ : io_requestor_2_req_bits_typ;
  assign io_mem_req_bits_cmd = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : T9;
  assign T9 = io_requestor_1_req_valid ? io_requestor_1_req_bits_cmd : io_requestor_2_req_bits_cmd;
  assign io_mem_req_bits_tag = T53;
  assign T53 = T10[4'h9:1'h0];
  assign T10 = io_requestor_0_req_valid ? T14 : T11;
  assign T11 = io_requestor_1_req_valid ? T13 : T12;
  assign T12 = {io_requestor_2_req_bits_tag, 2'h2};
  assign T13 = {io_requestor_1_req_bits_tag, 2'h1};
  assign T14 = {io_requestor_0_req_bits_tag, 2'h0};
  assign io_mem_req_bits_addr = T15;
  assign T15 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : T16;
  assign T16 = io_requestor_1_req_valid ? io_requestor_1_req_bits_addr : io_requestor_2_req_bits_addr;
  assign io_mem_req_valid = T17;
  assign T17 = T18 | io_requestor_2_req_valid;
  assign T18 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T54;
  assign T54 = {2'h0, T19};
  assign T19 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_0_replay_next_valid = T20;
  assign T20 = io_mem_replay_next_valid & T21;
  assign T21 = T22 == 2'h0;
  assign T22 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_replay = T23;
  assign T23 = io_mem_resp_bits_replay & T24;
  assign T24 = T25 == 2'h0;
  assign T25 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_0_resp_bits_nack = T26;
  assign T26 = io_mem_resp_bits_nack & T24;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T55;
  assign T55 = {2'h0, T27};
  assign T27 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_valid = T28;
  assign T28 = io_mem_resp_valid & T24;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T56;
  assign T56 = {2'h0, T29};
  assign T29 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_1_replay_next_valid = T30;
  assign T30 = io_mem_replay_next_valid & T31;
  assign T31 = T32 == 2'h1;
  assign T32 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_replay = T33;
  assign T33 = io_mem_resp_bits_replay & T34;
  assign T34 = T35 == 2'h1;
  assign T35 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_1_resp_bits_nack = T36;
  assign T36 = io_mem_resp_bits_nack & T34;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T57;
  assign T57 = {2'h0, T37};
  assign T37 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_valid = T38;
  assign T38 = io_mem_resp_valid & T34;
  assign io_requestor_1_req_ready = T39;
  assign T39 = io_requestor_0_req_ready & T40;
  assign T40 = io_requestor_0_req_valid ^ 1'h1;
  assign io_requestor_2_ordered = io_mem_ordered;
  assign io_requestor_2_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_2_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_2_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_2_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_2_replay_next_bits = T58;
  assign T58 = {2'h0, T41};
  assign T41 = io_mem_replay_next_bits >> 2'h2;
  assign io_requestor_2_replay_next_valid = T42;
  assign T42 = io_mem_replay_next_valid & T43;
  assign T43 = T44 == 2'h2;
  assign T44 = io_mem_replay_next_bits[1'h1:1'h0];
  assign io_requestor_2_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_2_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_2_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_2_resp_bits_replay = T45;
  assign T45 = io_mem_resp_bits_replay & T46;
  assign T46 = T47 == 2'h2;
  assign T47 = io_mem_resp_bits_tag[1'h1:1'h0];
  assign io_requestor_2_resp_bits_nack = T48;
  assign T48 = io_mem_resp_bits_nack & T46;
  assign io_requestor_2_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_2_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_2_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_2_resp_bits_tag = T59;
  assign T59 = {2'h0, T49};
  assign T49 = io_mem_resp_bits_tag >> 2'h2;
  assign io_requestor_2_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_2_resp_valid = T50;
  assign T50 = io_mem_resp_valid & T46;
  assign io_requestor_2_req_ready = T51;
  assign T51 = io_requestor_1_req_ready & T52;
  assign T52 = io_requestor_1_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_1 <= io_requestor_1_req_valid;
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module FPUDecoder(
    input [31:0] io_inst,
    output[4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap12,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_div,
    output io_sigs_sqrt,
    output io_sigs_round,
    output io_sigs_wflags
);

  wire T0;
  wire T1;
  wire[31:0] T2;
  wire T3;
  wire T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire T9;
  wire[31:0] T10;
  wire T11;
  wire T12;
  wire[31:0] T13;
  wire T14;
  wire T15;
  wire[31:0] T16;
  wire T17;
  wire[31:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire[31:0] T29;
  wire T30;
  wire T31;
  wire[31:0] T32;
  wire T33;
  wire[31:0] T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire[31:0] T41;
  wire T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire[31:0] T46;
  wire T47;
  wire[31:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire[31:0] T56;
  wire T57;
  wire[31:0] T58;
  wire T59;
  wire T60;
  wire[31:0] T61;
  wire T62;
  wire T63;
  wire[31:0] T64;
  wire T65;
  wire[31:0] T66;
  wire[4:0] T67;
  wire[3:0] T68;
  wire[2:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire[31:0] T75;
  wire T76;
  wire T77;
  wire[31:0] T78;
  wire T79;
  wire[31:0] T80;
  wire T81;
  wire T82;
  wire[31:0] T83;
  wire T84;
  wire T85;
  wire[31:0] T86;
  wire T87;
  wire[31:0] T88;


  assign io_sigs_wflags = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 32'h80000000;
  assign T2 = io_inst & 32'hc0000004;
  assign T3 = T6 | T4;
  assign T4 = T5 == 32'h8000000;
  assign T5 = io_inst & 32'h8002000;
  assign T6 = T9 | T7;
  assign T7 = T8 == 32'h40;
  assign T8 = io_inst & 32'h50;
  assign T9 = T10 == 32'h0;
  assign T10 = io_inst & 32'h20000004;
  assign io_sigs_round = T11;
  assign T11 = T14 | T12;
  assign T12 = T13 == 32'h40000000;
  assign T13 = io_inst & 32'h40002000;
  assign T14 = T9 | T7;
  assign io_sigs_sqrt = T15;
  assign T15 = T16 == 32'h50000010;
  assign T16 = io_inst & 32'hd0000010;
  assign io_sigs_div = T17;
  assign T17 = T18 == 32'h18000010;
  assign T18 = io_inst & 32'h58000010;
  assign io_sigs_fma = T19;
  assign T19 = T20 | T7;
  assign T20 = T23 | T21;
  assign T21 = T22 == 32'h0;
  assign T22 = io_inst & 32'h68000004;
  assign T23 = T24 == 32'h0;
  assign T24 = io_inst & 32'h70000004;
  assign io_sigs_fastpipe = T25;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h40000010;
  assign T27 = io_inst & 32'hd0000010;
  assign T28 = T29 == 32'h20000010;
  assign T29 = io_inst & 32'ha0000010;
  assign io_sigs_toint = T30;
  assign T30 = T33 | T31;
  assign T31 = T32 == 32'h80000010;
  assign T32 = io_inst & 32'h90000010;
  assign T33 = T34 == 32'h20;
  assign T34 = io_inst & 32'h20;
  assign io_sigs_fromint = T35;
  assign T35 = T36 == 32'h90000010;
  assign T36 = io_inst & 32'h90000010;
  assign io_sigs_single = T37;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'h40;
  assign T39 = io_inst & 32'h2000040;
  assign T40 = T41 == 32'h0;
  assign T41 = io_inst & 32'h1040;
  assign io_sigs_swap23 = T42;
  assign T42 = T43 == 32'h10;
  assign T43 = io_inst & 32'h30000010;
  assign io_sigs_swap12 = T44;
  assign T44 = T47 | T45;
  assign T45 = T46 == 32'h50000010;
  assign T46 = io_inst & 32'h50000010;
  assign T47 = T48 == 32'h0;
  assign T48 = io_inst & 32'h40;
  assign io_sigs_ren3 = T7;
  assign io_sigs_ren2 = T49;
  assign T49 = T50 | T7;
  assign T50 = T51 | T33;
  assign T51 = T52 == 32'h0;
  assign T52 = io_inst & 32'h40000004;
  assign io_sigs_ren1 = T53;
  assign T53 = T54 | T7;
  assign T54 = T57 | T55;
  assign T55 = T56 == 32'h0;
  assign T56 = io_inst & 32'h10000004;
  assign T57 = T58 == 32'h0;
  assign T58 = io_inst & 32'h80000004;
  assign io_sigs_wen = T59;
  assign T59 = T62 | T60;
  assign T60 = T61 == 32'h10000000;
  assign T61 = io_inst & 32'h10000020;
  assign T62 = T65 | T63;
  assign T63 = T64 == 32'h0;
  assign T64 = io_inst & 32'h30;
  assign T65 = T66 == 32'h0;
  assign T66 = io_inst & 32'h80000020;
  assign io_sigs_ldst = T47;
  assign io_sigs_cmd = T67;
  assign T67 = {T87, T68};
  assign T68 = {T84, T69};
  assign T69 = {T81, T70};
  assign T70 = {T76, T71};
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h8000010;
  assign T73 = io_inst & 32'h8000010;
  assign T74 = T75 == 32'h4;
  assign T75 = io_inst & 32'h4;
  assign T76 = T79 | T77;
  assign T77 = T78 == 32'h10000010;
  assign T78 = io_inst & 32'h10000010;
  assign T79 = T80 == 32'h8;
  assign T80 = io_inst & 32'h8;
  assign T81 = T47 | T82;
  assign T82 = T83 == 32'h20000000;
  assign T83 = io_inst & 32'h20000000;
  assign T84 = T47 | T85;
  assign T85 = T86 == 32'h40000000;
  assign T86 = io_inst & 32'h40000000;
  assign T87 = T88 == 32'h0;
  assign T88 = io_inst & 32'h10;
endmodule

module MulAddRecFN_preMul_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[23:0] io_mulAddA,
    output[23:0] io_mulAddB,
    output[47:0] io_mulAddC,
    output[2:0] io_toPostMul_highExpA,
    output io_toPostMul_isNaN_isQuietNaNA,
    output[2:0] io_toPostMul_highExpB,
    output io_toPostMul_isNaN_isQuietNaNB,
    output io_toPostMul_signProd,
    output io_toPostMul_isZeroProd,
    output io_toPostMul_opSignC,
    output[2:0] io_toPostMul_highExpC,
    output io_toPostMul_isNaN_isQuietNaNC,
    output io_toPostMul_isCDominant,
    output io_toPostMul_CAlignDist_0,
    output[6:0] io_toPostMul_CAlignDist,
    output io_toPostMul_bit0AlignedNegSigC,
    output[25:0] io_toPostMul_highAlignedNegSigC,
    output[10:0] io_toPostMul_sExpSum,
    output[1:0] io_toPostMul_roundingMode
);

  wire[10:0] sExpSum;
  wire[10:0] sExpAlignedProd;
  wire[10:0] T0;
  wire[10:0] T1;
  wire[7:0] T2;
  wire[8:0] expB;
  wire[2:0] T3;
  wire[2:0] T92;
  wire T4;
  wire T5;
  wire[10:0] T93;
  wire[8:0] expA;
  wire[10:0] T94;
  wire[8:0] expC;
  wire CAlignDist_floor;
  wire T6;
  wire[10:0] sNatCAlignDist;
  wire[10:0] T95;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T7;
  wire isZeroA;
  wire[2:0] T8;
  wire[25:0] T9;
  wire[74:0] alignedNegSigC;
  wire[75:0] T10;
  wire T11;
  wire doSubMags;
  wire opSignC;
  wire T12;
  wire T13;
  wire signProd;
  wire T14;
  wire T15;
  wire signB;
  wire signA;
  wire T16;
  wire[23:0] T17;
  wire[23:0] CExtraMask;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[6:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[5:0] T25;
  wire[7:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[3:0] T29;
  wire[7:0] T30;
  wire[23:0] T31;
  wire[128:0] T32;
  wire[6:0] CAlignDist;
  wire[6:0] T33;
  wire[6:0] T34;
  wire T35;
  wire[9:0] T36;
  wire[7:0] T37;
  wire[7:0] T96;
  wire[3:0] T38;
  wire[7:0] T39;
  wire[7:0] T97;
  wire[5:0] T40;
  wire[7:0] T41;
  wire[7:0] T98;
  wire[6:0] T42;
  wire[15:0] T43;
  wire[15:0] T44;
  wire[15:0] T45;
  wire[14:0] T46;
  wire[15:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[13:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[11:0] T54;
  wire[15:0] T55;
  wire[15:0] T56;
  wire[15:0] T57;
  wire[7:0] T58;
  wire[15:0] T59;
  wire[15:0] T60;
  wire[15:0] T99;
  wire[7:0] T61;
  wire[15:0] T62;
  wire[15:0] T100;
  wire[11:0] T63;
  wire[15:0] T64;
  wire[15:0] T101;
  wire[13:0] T65;
  wire[15:0] T66;
  wire[15:0] T102;
  wire[14:0] T67;
  wire[23:0] sigC;
  wire[22:0] fractC;
  wire T68;
  wire isZeroC;
  wire[2:0] T69;
  wire[74:0] T70;
  wire[74:0] T71;
  wire[74:0] T72;
  wire[73:0] T73;
  wire[49:0] T74;
  wire[49:0] T103;
  wire[23:0] negSigC;
  wire[23:0] T75;
  wire T76;
  wire CAlignDist_0;
  wire T77;
  wire[9:0] T78;
  wire isCDominant;
  wire T79;
  wire T80;
  wire[9:0] T81;
  wire T82;
  wire T83;
  wire[2:0] T84;
  wire T85;
  wire[22:0] fractB;
  wire[2:0] T86;
  wire T87;
  wire[22:0] fractA;
  wire[2:0] T88;
  wire[47:0] T89;
  wire[23:0] sigB;
  wire T90;
  wire[23:0] sigA;
  wire T91;


  assign io_toPostMul_roundingMode = io_roundingMode;
  assign io_toPostMul_sExpSum = sExpSum;
  assign sExpSum = CAlignDist_floor ? T94 : sExpAlignedProd;
  assign sExpAlignedProd = T0 + 11'h1b;
  assign T0 = T93 + T1;
  assign T1 = {T3, T2};
  assign T2 = expB[3'h7:1'h0];
  assign expB = io_b[5'h1f:5'h17];
  assign T3 = 3'h0 - T92;
  assign T92 = {2'h0, T4};
  assign T4 = T5 ^ 1'h1;
  assign T5 = expB[4'h8];
  assign T93 = {2'h0, expA};
  assign expA = io_a[5'h1f:5'h17];
  assign T94 = {2'h0, expC};
  assign expC = io_c[5'h1f:5'h17];
  assign CAlignDist_floor = isZeroProd | T6;
  assign T6 = sNatCAlignDist[4'ha];
  assign sNatCAlignDist = sExpAlignedProd - T95;
  assign T95 = {2'h0, expC};
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T7 == 3'h0;
  assign T7 = expB[4'h8:3'h6];
  assign isZeroA = T8 == 3'h0;
  assign T8 = expA[4'h8:3'h6];
  assign io_toPostMul_highAlignedNegSigC = T9;
  assign T9 = alignedNegSigC[7'h4a:6'h31];
  assign alignedNegSigC = T10[7'h4a:1'h0];
  assign T10 = {T70, T11};
  assign T11 = T16 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T13 ^ T12;
  assign T12 = io_op[1'h0];
  assign T13 = io_c[6'h20];
  assign signProd = T15 ^ T14;
  assign T14 = io_op[1'h1];
  assign T15 = signA ^ signB;
  assign signB = io_b[6'h20];
  assign signA = io_a[6'h20];
  assign T16 = T17 != 24'h0;
  assign T17 = sigC & CExtraMask;
  assign CExtraMask = {T43, T18};
  assign T18 = T41 | T19;
  assign T19 = T20 & 8'haa;
  assign T20 = T21 << 1'h1;
  assign T21 = T22[3'h6:1'h0];
  assign T22 = T39 | T23;
  assign T23 = T24 & 8'hcc;
  assign T24 = T25 << 2'h2;
  assign T25 = T26[3'h5:1'h0];
  assign T26 = T37 | T27;
  assign T27 = T28 & 8'hf0;
  assign T28 = T29 << 3'h4;
  assign T29 = T30[2'h3:1'h0];
  assign T30 = T31[5'h17:5'h10];
  assign T31 = T32[7'h4d:6'h36];
  assign T32 = $signed(129'h100000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = CAlignDist_floor ? 7'h0 : T33;
  assign T33 = T35 ? T34 : 7'h4a;
  assign T34 = sNatCAlignDist[3'h6:1'h0];
  assign T35 = T36 < 10'h4a;
  assign T36 = sNatCAlignDist[4'h9:1'h0];
  assign T37 = T96 & 8'hf;
  assign T96 = {4'h0, T38};
  assign T38 = T30 >> 3'h4;
  assign T39 = T97 & 8'h33;
  assign T97 = {2'h0, T40};
  assign T40 = T26 >> 2'h2;
  assign T41 = T98 & 8'h55;
  assign T98 = {1'h0, T42};
  assign T42 = T22 >> 1'h1;
  assign T43 = T66 | T44;
  assign T44 = T45 & 16'haaaa;
  assign T45 = T46 << 1'h1;
  assign T46 = T47[4'he:1'h0];
  assign T47 = T64 | T48;
  assign T48 = T49 & 16'hcccc;
  assign T49 = T50 << 2'h2;
  assign T50 = T51[4'hd:1'h0];
  assign T51 = T62 | T52;
  assign T52 = T53 & 16'hf0f0;
  assign T53 = T54 << 3'h4;
  assign T54 = T55[4'hb:1'h0];
  assign T55 = T60 | T56;
  assign T56 = T57 & 16'hff00;
  assign T57 = T58 << 4'h8;
  assign T58 = T59[3'h7:1'h0];
  assign T59 = T31[4'hf:1'h0];
  assign T60 = T99 & 16'hff;
  assign T99 = {8'h0, T61};
  assign T61 = T59 >> 4'h8;
  assign T62 = T100 & 16'hf0f;
  assign T100 = {4'h0, T63};
  assign T63 = T55 >> 3'h4;
  assign T64 = T101 & 16'h3333;
  assign T101 = {2'h0, T65};
  assign T65 = T51 >> 2'h2;
  assign T66 = T102 & 16'h5555;
  assign T102 = {1'h0, T67};
  assign T67 = T47 >> 1'h1;
  assign sigC = {T68, fractC};
  assign fractC = io_c[5'h16:1'h0];
  assign T68 = isZeroC ^ 1'h1;
  assign isZeroC = T69 == 3'h0;
  assign T69 = expC[4'h8:3'h6];
  assign T70 = $signed(T71) >>> CAlignDist;
  assign T71 = T72;
  assign T72 = {doSubMags, T73};
  assign T73 = {negSigC, T74};
  assign T74 = 50'h0 - T103;
  assign T103 = {49'h0, doSubMags};
  assign negSigC = doSubMags ? T75 : sigC;
  assign T75 = ~ sigC;
  assign io_toPostMul_bit0AlignedNegSigC = T76;
  assign T76 = alignedNegSigC[1'h0];
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign CAlignDist_0 = CAlignDist_floor | T77;
  assign T77 = T78 == 10'h0;
  assign T78 = sNatCAlignDist[4'h9:1'h0];
  assign io_toPostMul_isCDominant = isCDominant;
  assign isCDominant = T82 & T79;
  assign T79 = CAlignDist_floor | T80;
  assign T80 = T81 < 10'h19;
  assign T81 = sNatCAlignDist[4'h9:1'h0];
  assign T82 = isZeroC ^ 1'h1;
  assign io_toPostMul_isNaN_isQuietNaNC = T83;
  assign T83 = fractC[5'h16];
  assign io_toPostMul_highExpC = T84;
  assign T84 = expC[4'h8:3'h6];
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isNaN_isQuietNaNB = T85;
  assign T85 = fractB[5'h16];
  assign fractB = io_b[5'h16:1'h0];
  assign io_toPostMul_highExpB = T86;
  assign T86 = expB[4'h8:3'h6];
  assign io_toPostMul_isNaN_isQuietNaNA = T87;
  assign T87 = fractA[5'h16];
  assign fractA = io_a[5'h16:1'h0];
  assign io_toPostMul_highExpA = T88;
  assign T88 = expA[4'h8:3'h6];
  assign io_mulAddC = T89;
  assign T89 = alignedNegSigC[6'h30:1'h1];
  assign io_mulAddB = sigB;
  assign sigB = {T90, fractB};
  assign T90 = isZeroB ^ 1'h1;
  assign io_mulAddA = sigA;
  assign sigA = {T91, fractA};
  assign T91 = isZeroA ^ 1'h1;
endmodule

module MulAddRecFN_postMul_0(
    input [2:0] io_fromPreMul_highExpA,
    input  io_fromPreMul_isNaN_isQuietNaNA,
    input [2:0] io_fromPreMul_highExpB,
    input  io_fromPreMul_isNaN_isQuietNaNB,
    input  io_fromPreMul_signProd,
    input  io_fromPreMul_isZeroProd,
    input  io_fromPreMul_opSignC,
    input [2:0] io_fromPreMul_highExpC,
    input  io_fromPreMul_isNaN_isQuietNaNC,
    input  io_fromPreMul_isCDominant,
    input  io_fromPreMul_CAlignDist_0,
    input [6:0] io_fromPreMul_CAlignDist,
    input  io_fromPreMul_bit0AlignedNegSigC,
    input [25:0] io_fromPreMul_highAlignedNegSigC,
    input [10:0] io_fromPreMul_sExpSum,
    input [1:0] io_fromPreMul_roundingMode,
    input [48:0] io_mulAddResult,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[27:0] T4;
  wire[27:0] T359;
  wire[25:0] T5;
  wire[26:0] roundMask;
  wire[26:0] T6;
  wire[24:0] T7;
  wire[24:0] T360;
  wire T8;
  wire[24:0] T9;
  wire[8:0] T10;
  wire T11;
  wire[8:0] T12;
  wire[24:0] T13;
  wire[1024:0] T14;
  wire[9:0] T15;
  wire[9:0] sExpX3_13;
  wire[10:0] sExpX3;
  wire[10:0] T361;
  wire[6:0] estNormDist;
  wire[6:0] T16;
  wire[6:0] estNormNeg_dist;
  wire[6:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[5:0] T365;
  wire[5:0] T366;
  wire[5:0] T367;
  wire[5:0] T368;
  wire[5:0] T369;
  wire[5:0] T370;
  wire[5:0] T371;
  wire[5:0] T372;
  wire[5:0] T373;
  wire[5:0] T374;
  wire[5:0] T375;
  wire[5:0] T376;
  wire[5:0] T377;
  wire[5:0] T378;
  wire[5:0] T379;
  wire[5:0] T380;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire[4:0] T385;
  wire[4:0] T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire[4:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[4:0] T392;
  wire[4:0] T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire[4:0] T396;
  wire[3:0] T397;
  wire[3:0] T398;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[2:0] T405;
  wire[2:0] T406;
  wire[2:0] T407;
  wire[2:0] T408;
  wire[1:0] T409;
  wire[1:0] T410;
  wire T411;
  wire[49:0] T18;
  wire[49:0] T19;
  wire[50:0] T20;
  wire[50:0] T21;
  wire[49:0] T22;
  wire[49:0] T23;
  wire[74:0] sigSum;
  wire[48:0] T24;
  wire[47:0] T25;
  wire[25:0] T26;
  wire[25:0] T27;
  wire T28;
  wire[50:0] T412;
  wire[49:0] T29;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire notCDom_signSigSum;
  wire[6:0] CDom_estNormDist;
  wire[6:0] T461;
  wire[4:0] T30;
  wire[6:0] T31;
  wire T32;
  wire doSubMags;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[6:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[5:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[3:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[7:0] T462;
  wire[3:0] T47;
  wire[7:0] T48;
  wire[7:0] T463;
  wire[5:0] T49;
  wire[7:0] T50;
  wire[7:0] T464;
  wire[6:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[15:0] T54;
  wire[14:0] T55;
  wire[15:0] T56;
  wire[15:0] T57;
  wire[15:0] T58;
  wire[13:0] T59;
  wire[15:0] T60;
  wire[15:0] T61;
  wire[15:0] T62;
  wire[11:0] T63;
  wire[15:0] T64;
  wire[15:0] T65;
  wire[15:0] T66;
  wire[7:0] T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire[15:0] T465;
  wire[7:0] T70;
  wire[15:0] T71;
  wire[15:0] T466;
  wire[11:0] T72;
  wire[15:0] T73;
  wire[15:0] T467;
  wire[13:0] T74;
  wire[15:0] T75;
  wire[15:0] T468;
  wire[14:0] T76;
  wire[26:0] T77;
  wire[26:0] T469;
  wire T78;
  wire[27:0] sigX3;
  wire[42:0] T79;
  wire T80;
  wire T81;
  wire[15:0] T82;
  wire[15:0] absSigSumExtraMask;
  wire[14:0] T83;
  wire[6:0] T84;
  wire[2:0] T85;
  wire T86;
  wire[2:0] T87;
  wire[6:0] T88;
  wire[14:0] T89;
  wire[16:0] T90;
  wire[3:0] normTo2ShiftDist;
  wire[3:0] estNormDist_5;
  wire[1:0] T91;
  wire T92;
  wire[1:0] T93;
  wire T94;
  wire[3:0] T95;
  wire[1:0] T96;
  wire T97;
  wire[1:0] T98;
  wire[3:0] T99;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire[1:0] T103;
  wire T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[6:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[5:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[3:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T470;
  wire[3:0] T119;
  wire[7:0] T120;
  wire[7:0] T471;
  wire[5:0] T121;
  wire[7:0] T122;
  wire[7:0] T472;
  wire[6:0] T123;
  wire[15:0] T124;
  wire[42:0] cFirstNormAbsSigSum;
  wire[42:0] T473;
  wire[41:0] T125;
  wire[41:0] notCDom_pos_firstNormAbsSigSum;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[31:0] T128;
  wire[31:0] T474;
  wire[9:0] T129;
  wire[41:0] T475;
  wire[33:0] T130;
  wire T131;
  wire T132;
  wire[1:0] firstReduceSigSum;
  wire T133;
  wire[17:0] T134;
  wire T135;
  wire[15:0] T136;
  wire T137;
  wire T138;
  wire[1:0] firstReduceComplSigSum;
  wire T139;
  wire[17:0] T140;
  wire[74:0] complSigSum;
  wire T141;
  wire[15:0] T142;
  wire[32:0] T143;
  wire T144;
  wire[41:0] T145;
  wire[41:0] T146;
  wire[41:0] T147;
  wire[15:0] T148;
  wire[15:0] T476;
  wire[25:0] T149;
  wire T150;
  wire T151;
  wire[41:0] CDom_firstNormAbsSigSum;
  wire[41:0] T152;
  wire[41:0] T153;
  wire T154;
  wire[40:0] T155;
  wire T156;
  wire T157;
  wire[41:0] T158;
  wire[41:0] T159;
  wire[41:0] T160;
  wire T161;
  wire[40:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire[41:0] T166;
  wire[41:0] T167;
  wire[41:0] T168;
  wire T169;
  wire[40:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire[41:0] T174;
  wire[41:0] T175;
  wire T176;
  wire[40:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[42:0] T182;
  wire[42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[42:0] T183;
  wire[42:0] T184;
  wire[10:0] T185;
  wire[42:0] T477;
  wire[32:0] T186;
  wire T187;
  wire[31:0] T188;
  wire T189;
  wire[42:0] T190;
  wire[42:0] T478;
  wire[41:0] T191;
  wire[42:0] T192;
  wire[26:0] T193;
  wire T194;
  wire T195;
  wire[42:0] T479;
  wire T196;
  wire[15:0] T197;
  wire[15:0] T198;
  wire[15:0] T199;
  wire[41:0] T200;
  wire[41:0] T201;
  wire roundPosBit;
  wire[27:0] T202;
  wire[27:0] T480;
  wire[26:0] roundPosMask;
  wire[26:0] T481;
  wire[25:0] T203;
  wire[25:0] T204;
  wire T205;
  wire allRound;
  wire allRoundExtra;
  wire[27:0] T206;
  wire[27:0] T482;
  wire[25:0] T207;
  wire[27:0] T208;
  wire doIncrSig;
  wire T209;
  wire T210;
  wire T211;
  wire commonCase;
  wire T212;
  wire notSpecial_addZeros;
  wire isZeroC;
  wire T213;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T214;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T215;
  wire isSpecialA;
  wire[1:0] T216;
  wire underflow;
  wire underflowY;
  wire T217;
  wire T218;
  wire[9:0] T483;
  wire[7:0] T219;
  wire sigX3Shift1;
  wire[1:0] T220;
  wire T221;
  wire overflow;
  wire overflowY;
  wire[2:0] T222;
  wire[10:0] sExpY;
  wire[10:0] T223;
  wire[10:0] T224;
  wire T225;
  wire[1:0] T226;
  wire[25:0] sigY3;
  wire[25:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[25:0] T230;
  wire[25:0] roundUp_sigY3;
  wire[25:0] T231;
  wire[25:0] T232;
  wire[27:0] T233;
  wire[27:0] T484;
  wire roundEven;
  wire T234;
  wire T235;
  wire T236;
  wire roundingMode_nearest_even;
  wire T237;
  wire T238;
  wire T239;
  wire[25:0] T240;
  wire[25:0] T241;
  wire roundUp;
  wire T242;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T243;
  wire doNegSignSum;
  wire T244;
  wire T245;
  wire isZeroY;
  wire[2:0] T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[25:0] T260;
  wire[25:0] T261;
  wire[27:0] T262;
  wire[27:0] T485;
  wire[26:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[10:0] T267;
  wire[10:0] T268;
  wire T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire[1:0] T273;
  wire invalid;
  wire notSigNaN_invalid;
  wire T274;
  wire T275;
  wire isInfC;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire isInfB;
  wire T280;
  wire T281;
  wire isInfA;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire isNaNB;
  wire T286;
  wire T287;
  wire isNaNA;
  wire T288;
  wire T289;
  wire T290;
  wire isZeroA;
  wire T291;
  wire isZeroB;
  wire T292;
  wire isSigNaNC;
  wire T293;
  wire isNaNC;
  wire T294;
  wire T295;
  wire isSigNaNB;
  wire T296;
  wire isSigNaNA;
  wire T297;
  wire[32:0] T298;
  wire[31:0] T299;
  wire[22:0] fractOut;
  wire[22:0] T300;
  wire[22:0] T486;
  wire pegMaxFiniteMagOut;
  wire T301;
  wire overflowY_roundMagUp;
  wire roundMagUp;
  wire T302;
  wire T303;
  wire T304;
  wire[22:0] T305;
  wire[22:0] fractY;
  wire[22:0] T306;
  wire[22:0] T307;
  wire[22:0] T308;
  wire isNaNOut;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire totalUnderflowY;
  wire T313;
  wire T314;
  wire[8:0] T315;
  wire T316;
  wire T317;
  wire[8:0] expOut;
  wire[8:0] T318;
  wire[8:0] T319;
  wire[8:0] T320;
  wire notNaN_isInfOut;
  wire T321;
  wire T322;
  wire T323;
  wire[8:0] T324;
  wire[8:0] T325;
  wire[8:0] T326;
  wire[8:0] T327;
  wire pegMinFiniteMagOut;
  wire T328;
  wire[8:0] T329;
  wire[8:0] T330;
  wire[8:0] T331;
  wire[8:0] T332;
  wire[8:0] T333;
  wire[8:0] T334;
  wire[8:0] T335;
  wire[8:0] T336;
  wire[8:0] T337;
  wire[8:0] T338;
  wire[8:0] T339;
  wire[8:0] T340;
  wire notSpecial_isZeroOut;
  wire T341;
  wire[8:0] expY;
  wire signOut;
  wire T342;
  wire T343;
  wire uncommonCaseSignOut;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;


  assign io_exceptionFlags = T0;
  assign T0 = {T273, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T205 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 28'h0;
  assign T4 = sigX3 & T359;
  assign T359 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T77 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T360;
  assign T360 = {24'h0, T8};
  assign T8 = sigX3[5'h1a];
  assign T9 = {T52, T10};
  assign T10 = {T33, T11};
  assign T11 = T12[4'h8];
  assign T12 = T13[5'h18:5'h10];
  assign T13 = T14[8'h83:7'h6b];
  assign T14 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T15;
  assign T15 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'h9:1'h0];
  assign sExpX3 = io_fromPreMul_sExpSum - T361;
  assign T361 = {4'h0, estNormDist};
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : T16;
  assign T16 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = 7'h49 - T362;
  assign T362 = {1'h0, T363};
  assign T363 = T460 ? 6'h31 : T364;
  assign T364 = T459 ? 6'h30 : T365;
  assign T365 = T458 ? 6'h2f : T366;
  assign T366 = T457 ? 6'h2e : T367;
  assign T367 = T456 ? 6'h2d : T368;
  assign T368 = T455 ? 6'h2c : T369;
  assign T369 = T454 ? 6'h2b : T370;
  assign T370 = T453 ? 6'h2a : T371;
  assign T371 = T452 ? 6'h29 : T372;
  assign T372 = T451 ? 6'h28 : T373;
  assign T373 = T450 ? 6'h27 : T374;
  assign T374 = T449 ? 6'h26 : T375;
  assign T375 = T448 ? 6'h25 : T376;
  assign T376 = T447 ? 6'h24 : T377;
  assign T377 = T446 ? 6'h23 : T378;
  assign T378 = T445 ? 6'h22 : T379;
  assign T379 = T444 ? 6'h21 : T380;
  assign T380 = T443 ? 6'h20 : T381;
  assign T381 = T442 ? 5'h1f : T382;
  assign T382 = T441 ? 5'h1e : T383;
  assign T383 = T440 ? 5'h1d : T384;
  assign T384 = T439 ? 5'h1c : T385;
  assign T385 = T438 ? 5'h1b : T386;
  assign T386 = T437 ? 5'h1a : T387;
  assign T387 = T436 ? 5'h19 : T388;
  assign T388 = T435 ? 5'h18 : T389;
  assign T389 = T434 ? 5'h17 : T390;
  assign T390 = T433 ? 5'h16 : T391;
  assign T391 = T432 ? 5'h15 : T392;
  assign T392 = T431 ? 5'h14 : T393;
  assign T393 = T430 ? 5'h13 : T394;
  assign T394 = T429 ? 5'h12 : T395;
  assign T395 = T428 ? 5'h11 : T396;
  assign T396 = T427 ? 5'h10 : T397;
  assign T397 = T426 ? 4'hf : T398;
  assign T398 = T425 ? 4'he : T399;
  assign T399 = T424 ? 4'hd : T400;
  assign T400 = T423 ? 4'hc : T401;
  assign T401 = T422 ? 4'hb : T402;
  assign T402 = T421 ? 4'ha : T403;
  assign T403 = T420 ? 4'h9 : T404;
  assign T404 = T419 ? 4'h8 : T405;
  assign T405 = T418 ? 3'h7 : T406;
  assign T406 = T417 ? 3'h6 : T407;
  assign T407 = T416 ? 3'h5 : T408;
  assign T408 = T415 ? 3'h4 : T409;
  assign T409 = T414 ? 2'h3 : T410;
  assign T410 = T413 ? 2'h2 : T411;
  assign T411 = T18[1'h1];
  assign T18 = T19;
  assign T19 = T20[6'h31:1'h0];
  assign T20 = T412 ^ T21;
  assign T21 = T22 << 1'h1;
  assign T22 = 50'h0 | T23;
  assign T23 = sigSum[6'h32:1'h1];
  assign sigSum = {T26, T24};
  assign T24 = {T25, io_fromPreMul_bit0AlignedNegSigC};
  assign T25 = io_mulAddResult[6'h2f:1'h0];
  assign T26 = T28 ? T27 : io_fromPreMul_highAlignedNegSigC;
  assign T27 = io_fromPreMul_highAlignedNegSigC + 26'h1;
  assign T28 = io_mulAddResult[6'h30];
  assign T412 = {1'h0, T29};
  assign T29 = 50'h0 ^ T23;
  assign T413 = T18[2'h2];
  assign T414 = T18[2'h3];
  assign T415 = T18[3'h4];
  assign T416 = T18[3'h5];
  assign T417 = T18[3'h6];
  assign T418 = T18[3'h7];
  assign T419 = T18[4'h8];
  assign T420 = T18[4'h9];
  assign T421 = T18[4'ha];
  assign T422 = T18[4'hb];
  assign T423 = T18[4'hc];
  assign T424 = T18[4'hd];
  assign T425 = T18[4'he];
  assign T426 = T18[4'hf];
  assign T427 = T18[5'h10];
  assign T428 = T18[5'h11];
  assign T429 = T18[5'h12];
  assign T430 = T18[5'h13];
  assign T431 = T18[5'h14];
  assign T432 = T18[5'h15];
  assign T433 = T18[5'h16];
  assign T434 = T18[5'h17];
  assign T435 = T18[5'h18];
  assign T436 = T18[5'h19];
  assign T437 = T18[5'h1a];
  assign T438 = T18[5'h1b];
  assign T439 = T18[5'h1c];
  assign T440 = T18[5'h1d];
  assign T441 = T18[5'h1e];
  assign T442 = T18[5'h1f];
  assign T443 = T18[6'h20];
  assign T444 = T18[6'h21];
  assign T445 = T18[6'h22];
  assign T446 = T18[6'h23];
  assign T447 = T18[6'h24];
  assign T448 = T18[6'h25];
  assign T449 = T18[6'h26];
  assign T450 = T18[6'h27];
  assign T451 = T18[6'h28];
  assign T452 = T18[6'h29];
  assign T453 = T18[6'h2a];
  assign T454 = T18[6'h2b];
  assign T455 = T18[6'h2c];
  assign T456 = T18[6'h2d];
  assign T457 = T18[6'h2e];
  assign T458 = T18[6'h2f];
  assign T459 = T18[6'h30];
  assign T460 = T18[6'h31];
  assign notCDom_signSigSum = sigSum[6'h33];
  assign CDom_estNormDist = T32 ? io_fromPreMul_CAlignDist : T461;
  assign T461 = {2'h0, T30};
  assign T30 = T31[3'h4:1'h0];
  assign T31 = io_fromPreMul_CAlignDist - 7'h1;
  assign T32 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T33 = T50 | T34;
  assign T34 = T35 & 8'haa;
  assign T35 = T36 << 1'h1;
  assign T36 = T37[3'h6:1'h0];
  assign T37 = T48 | T38;
  assign T38 = T39 & 8'hcc;
  assign T39 = T40 << 2'h2;
  assign T40 = T41[3'h5:1'h0];
  assign T41 = T46 | T42;
  assign T42 = T43 & 8'hf0;
  assign T43 = T44 << 3'h4;
  assign T44 = T45[2'h3:1'h0];
  assign T45 = T12[3'h7:1'h0];
  assign T46 = T462 & 8'hf;
  assign T462 = {4'h0, T47};
  assign T47 = T45 >> 3'h4;
  assign T48 = T463 & 8'h33;
  assign T463 = {2'h0, T49};
  assign T49 = T41 >> 2'h2;
  assign T50 = T464 & 8'h55;
  assign T464 = {1'h0, T51};
  assign T51 = T37 >> 1'h1;
  assign T52 = T75 | T53;
  assign T53 = T54 & 16'haaaa;
  assign T54 = T55 << 1'h1;
  assign T55 = T56[4'he:1'h0];
  assign T56 = T73 | T57;
  assign T57 = T58 & 16'hcccc;
  assign T58 = T59 << 2'h2;
  assign T59 = T60[4'hd:1'h0];
  assign T60 = T71 | T61;
  assign T61 = T62 & 16'hf0f0;
  assign T62 = T63 << 3'h4;
  assign T63 = T64[4'hb:1'h0];
  assign T64 = T69 | T65;
  assign T65 = T66 & 16'hff00;
  assign T66 = T67 << 4'h8;
  assign T67 = T68[3'h7:1'h0];
  assign T68 = T13[4'hf:1'h0];
  assign T69 = T465 & 16'hff;
  assign T465 = {8'h0, T70};
  assign T70 = T68 >> 4'h8;
  assign T71 = T466 & 16'hf0f;
  assign T466 = {4'h0, T72};
  assign T72 = T64 >> 3'h4;
  assign T73 = T467 & 16'h3333;
  assign T467 = {2'h0, T74};
  assign T74 = T60 >> 2'h2;
  assign T75 = T468 & 16'h5555;
  assign T468 = {1'h0, T76};
  assign T76 = T56 >> 1'h1;
  assign T77 = 27'h0 - T469;
  assign T469 = {26'h0, T78};
  assign T78 = sExpX3[4'ha];
  assign sigX3 = T79[5'h1b:1'h0];
  assign T79 = {T200, T80};
  assign T80 = doIncrSig ? T196 : T81;
  assign T81 = T82 != 16'h0;
  assign T82 = T124 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T83, 1'h1};
  assign T83 = {T105, T84};
  assign T84 = {T95, T85};
  assign T85 = {T91, T86};
  assign T86 = T87[2'h2];
  assign T87 = T88[3'h6:3'h4];
  assign T88 = T89[4'he:4'h8];
  assign T89 = T90[4'hf:1'h1];
  assign T90 = $signed(17'h10000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = estNormDist[2'h3:1'h0];
  assign T91 = {T94, T92};
  assign T92 = T93[1'h1];
  assign T93 = T87[1'h1:1'h0];
  assign T94 = T93[1'h0];
  assign T95 = {T101, T96};
  assign T96 = {T100, T97};
  assign T97 = T98[1'h1];
  assign T98 = T99[2'h3:2'h2];
  assign T99 = T88[2'h3:1'h0];
  assign T100 = T98[1'h0];
  assign T101 = {T104, T102};
  assign T102 = T103[1'h1];
  assign T103 = T99[1'h1:1'h0];
  assign T104 = T103[1'h0];
  assign T105 = T122 | T106;
  assign T106 = T107 & 8'haa;
  assign T107 = T108 << 1'h1;
  assign T108 = T109[3'h6:1'h0];
  assign T109 = T120 | T110;
  assign T110 = T111 & 8'hcc;
  assign T111 = T112 << 2'h2;
  assign T112 = T113[3'h5:1'h0];
  assign T113 = T118 | T114;
  assign T114 = T115 & 8'hf0;
  assign T115 = T116 << 3'h4;
  assign T116 = T117[2'h3:1'h0];
  assign T117 = T89[3'h7:1'h0];
  assign T118 = T470 & 8'hf;
  assign T470 = {4'h0, T119};
  assign T119 = T117 >> 3'h4;
  assign T120 = T471 & 8'h33;
  assign T471 = {2'h0, T121};
  assign T121 = T113 >> 2'h2;
  assign T122 = T472 & 8'h55;
  assign T472 = {1'h0, T123};
  assign T123 = T109 >> 1'h1;
  assign T124 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T182 : T473;
  assign T473 = {1'h0, T125};
  assign T125 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T151 ? T145 : T126;
  assign T126 = T144 ? T475 : T127;
  assign T127 = {T129, T128};
  assign T128 = 32'h0 - T474;
  assign T474 = {31'h0, doSubMags};
  assign T129 = sigSum[4'ha:1'h1];
  assign T475 = {8'h0, T130};
  assign T130 = {T143, T131};
  assign T131 = doSubMags ? T137 : T132;
  assign T132 = firstReduceSigSum[1'h0];
  assign firstReduceSigSum = {T135, T133};
  assign T133 = T134 != 18'h0;
  assign T134 = sigSum[5'h11:1'h0];
  assign T135 = T136 != 16'h0;
  assign T136 = sigSum[6'h21:5'h12];
  assign T137 = T138 ^ 1'h1;
  assign T138 = firstReduceComplSigSum[1'h0];
  assign firstReduceComplSigSum = {T141, T139};
  assign T139 = T140 != 18'h0;
  assign T140 = complSigSum[5'h11:1'h0];
  assign complSigSum = ~ sigSum;
  assign T141 = T142 != 16'h0;
  assign T142 = complSigSum[6'h21:5'h12];
  assign T143 = sigSum[6'h32:5'h12];
  assign T144 = estNormNeg_dist[3'h4];
  assign T145 = T150 ? T147 : T146;
  assign T146 = sigSum[6'h2a:1'h1];
  assign T147 = {T149, T148};
  assign T148 = 16'h0 - T476;
  assign T476 = {15'h0, doSubMags};
  assign T149 = sigSum[5'h1a:1'h1];
  assign T150 = estNormNeg_dist[3'h4];
  assign T151 = estNormNeg_dist[3'h5];
  assign CDom_firstNormAbsSigSum = T158 | T152;
  assign T152 = T156 ? T153 : 42'h0;
  assign T153 = {T155, T154};
  assign T154 = firstReduceComplSigSum[1'h0];
  assign T155 = complSigSum[6'h3a:5'h12];
  assign T156 = doSubMags & T157;
  assign T157 = CDom_estNormDist[3'h4];
  assign T158 = T166 | T159;
  assign T159 = T163 ? T160 : 42'h0;
  assign T160 = {T162, T161};
  assign T161 = firstReduceComplSigSum != 2'h0;
  assign T162 = complSigSum[7'h4a:6'h22];
  assign T163 = doSubMags & T164;
  assign T164 = T165 ^ 1'h1;
  assign T165 = CDom_estNormDist[3'h4];
  assign T166 = T174 | T167;
  assign T167 = T171 ? T168 : 42'h0;
  assign T168 = {T170, T169};
  assign T169 = firstReduceSigSum[1'h0];
  assign T170 = sigSum[6'h3a:5'h12];
  assign T171 = T173 & T172;
  assign T172 = CDom_estNormDist[3'h4];
  assign T173 = doSubMags ^ 1'h1;
  assign T174 = T178 ? T175 : 42'h0;
  assign T175 = {T177, T176};
  assign T176 = firstReduceSigSum != 2'h0;
  assign T177 = sigSum[7'h4a:6'h22];
  assign T178 = T181 & T179;
  assign T179 = T180 ^ 1'h1;
  assign T180 = CDom_estNormDist[3'h4];
  assign T181 = doSubMags ^ 1'h1;
  assign T182 = io_fromPreMul_isCDominant ? T479 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T195 ? T190 : T183;
  assign T183 = T189 ? T477 : T184;
  assign T184 = T185 << 6'h20;
  assign T185 = complSigSum[4'hb:1'h1];
  assign T477 = {10'h0, T186};
  assign T186 = {T188, T187};
  assign T187 = firstReduceComplSigSum[1'h0];
  assign T188 = complSigSum[6'h31:5'h12];
  assign T189 = estNormNeg_dist[3'h4];
  assign T190 = T194 ? T192 : T478;
  assign T478 = {1'h0, T191};
  assign T191 = complSigSum[6'h2a:1'h1];
  assign T192 = T193 << 5'h10;
  assign T193 = complSigSum[5'h1b:1'h1];
  assign T194 = estNormNeg_dist[3'h4];
  assign T195 = estNormNeg_dist[3'h5];
  assign T479 = {1'h0, CDom_firstNormAbsSigSum};
  assign T196 = T197 == 16'h0;
  assign T197 = T198 & absSigSumExtraMask;
  assign T198 = ~ T199;
  assign T199 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign T200 = T201 >> normTo2ShiftDist;
  assign T201 = cFirstNormAbsSigSum[6'h2a:1'h1];
  assign roundPosBit = T202 != 28'h0;
  assign T202 = sigX3 & T480;
  assign T480 = {1'h0, roundPosMask};
  assign roundPosMask = T481 & roundMask;
  assign T481 = {1'h0, T203};
  assign T203 = ~ T204;
  assign T204 = roundMask >> 1'h1;
  assign T205 = allRound ^ 1'h1;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T206 == 28'h0;
  assign T206 = T208 & T482;
  assign T482 = {2'h0, T207};
  assign T207 = roundMask >> 1'h1;
  assign T208 = ~ sigX3;
  assign doIncrSig = T209 & doSubMags;
  assign T209 = T211 & T210;
  assign T210 = notCDom_signSigSum ^ 1'h1;
  assign T211 = io_fromPreMul_isCDominant ^ 1'h1;
  assign commonCase = T213 & T212;
  assign T212 = notSpecial_addZeros ^ 1'h1;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign isZeroC = io_fromPreMul_highExpC == 3'h0;
  assign T213 = addSpecial ^ 1'h1;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T214 == 2'h3;
  assign T214 = io_fromPreMul_highExpC[2'h2:1'h1];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T215 == 2'h3;
  assign T215 = io_fromPreMul_highExpB[2'h2:1'h1];
  assign isSpecialA = T216 == 2'h3;
  assign T216 = io_fromPreMul_highExpA[2'h2:1'h1];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T217;
  assign T217 = T221 | T218;
  assign T218 = sExpX3_13 <= T483;
  assign T483 = {2'h0, T219};
  assign T219 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign sigX3Shift1 = T220 == 2'h0;
  assign T220 = sigX3[5'h1b:5'h1a];
  assign T221 = sExpX3[4'ha];
  assign overflow = commonCase & overflowY;
  assign overflowY = T222 == 3'h3;
  assign T222 = sExpY[4'h9:3'h7];
  assign sExpY = T267 | T223;
  assign T223 = T225 ? T224 : 11'h0;
  assign T224 = sExpX3 - 11'h1;
  assign T225 = T226 == 2'h0;
  assign T226 = sigY3[5'h19:5'h18];
  assign sigY3 = T240 | T227;
  assign T227 = roundEven ? T228 : 26'h0;
  assign T228 = roundUp_sigY3 & T229;
  assign T229 = ~ T230;
  assign T230 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T231;
  assign T231 = T232 + 26'h1;
  assign T232 = T233 >> 2'h2;
  assign T233 = sigX3 | T484;
  assign T484 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T237 : T234;
  assign T234 = T236 & T235;
  assign T235 = anyRoundExtra ^ 1'h1;
  assign T236 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign T237 = T238 & allRoundExtra;
  assign T238 = roundingMode_nearest_even & T239;
  assign T239 = roundPosBit ^ 1'h1;
  assign T240 = T260 | T241;
  assign T241 = roundUp ? roundUp_sigY3 : 26'h0;
  assign roundUp = T247 | T242;
  assign T242 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign signY = isZeroY ? roundingMode_min : T243;
  assign T243 = io_fromPreMul_signProd ^ doNegSignSum;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T244 : notCDom_signSigSum;
  assign T244 = doSubMags & T245;
  assign T245 = isZeroC ^ 1'h1;
  assign isZeroY = T246 == 3'h0;
  assign T246 = sigX3[5'h1b:5'h19];
  assign T247 = T250 | T248;
  assign T248 = T249 & roundPosBit;
  assign T249 = doIncrSig & roundingMode_nearest_even;
  assign T250 = T252 | T251;
  assign T251 = doIncrSig & allRound;
  assign T252 = T256 | T253;
  assign T253 = T254 & anyRound;
  assign T254 = T255 & roundDirectUp;
  assign T255 = doIncrSig ^ 1'h1;
  assign T256 = T257 & anyRoundExtra;
  assign T257 = T258 & roundPosBit;
  assign T258 = T259 & roundingMode_nearest_even;
  assign T259 = doIncrSig ^ 1'h1;
  assign T260 = T264 ? T261 : 26'h0;
  assign T261 = T262 >> 2'h2;
  assign T262 = sigX3 & T485;
  assign T485 = {1'h0, T263};
  assign T263 = ~ roundMask;
  assign T264 = T266 & T265;
  assign T265 = roundEven ^ 1'h1;
  assign T266 = roundUp ^ 1'h1;
  assign T267 = T270 | T268;
  assign T268 = T269 ? sExpX3 : 11'h0;
  assign T269 = sigY3[5'h18];
  assign T270 = T272 ? T271 : 11'h0;
  assign T271 = sExpX3 + 11'h1;
  assign T272 = sigY3[5'h19];
  assign T273 = {invalid, 1'h0};
  assign invalid = T292 | notSigNaN_invalid;
  assign notSigNaN_invalid = T289 | T274;
  assign T274 = T275 & doSubMags;
  assign T275 = T278 & isInfC;
  assign isInfC = isSpecialC & T276;
  assign T276 = T277 ^ 1'h1;
  assign T277 = io_fromPreMul_highExpC[1'h0];
  assign T278 = T284 & T279;
  assign T279 = isInfA | isInfB;
  assign isInfB = isSpecialB & T280;
  assign T280 = T281 ^ 1'h1;
  assign T281 = io_fromPreMul_highExpB[1'h0];
  assign isInfA = isSpecialA & T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = io_fromPreMul_highExpA[1'h0];
  assign T284 = T287 & T285;
  assign T285 = isNaNB ^ 1'h1;
  assign isNaNB = isSpecialB & T286;
  assign T286 = io_fromPreMul_highExpB[1'h0];
  assign T287 = isNaNA ^ 1'h1;
  assign isNaNA = isSpecialA & T288;
  assign T288 = io_fromPreMul_highExpA[1'h0];
  assign T289 = T291 | T290;
  assign T290 = isZeroA & isInfB;
  assign isZeroA = io_fromPreMul_highExpA == 3'h0;
  assign T291 = isInfA & isZeroB;
  assign isZeroB = io_fromPreMul_highExpB == 3'h0;
  assign T292 = T295 | isSigNaNC;
  assign isSigNaNC = isNaNC & T293;
  assign T293 = io_fromPreMul_isNaN_isQuietNaNC ^ 1'h1;
  assign isNaNC = isSpecialC & T294;
  assign T294 = io_fromPreMul_highExpC[1'h0];
  assign T295 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T296;
  assign T296 = io_fromPreMul_isNaN_isQuietNaNB ^ 1'h1;
  assign isSigNaNA = isNaNA & T297;
  assign T297 = io_fromPreMul_isNaN_isQuietNaNA ^ 1'h1;
  assign io_out = T298;
  assign T298 = {signOut, T299};
  assign T299 = {expOut, fractOut};
  assign fractOut = T305 | T300;
  assign T300 = 23'h0 - T486;
  assign T486 = {22'h0, pegMaxFiniteMagOut};
  assign pegMaxFiniteMagOut = overflow & T301;
  assign T301 = overflowY_roundMagUp ^ 1'h1;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign roundMagUp = T304 | T302;
  assign T302 = roundingMode_max & T303;
  assign T303 = signY ^ 1'h1;
  assign T304 = roundingMode_min & signY;
  assign T305 = T311 ? T308 : fractY;
  assign fractY = sigX3Shift1 ? T307 : T306;
  assign T306 = sigY3[5'h17:1'h1];
  assign T307 = sigY3[5'h16:1'h0];
  assign T308 = isNaNOut ? 23'h400000 : 23'h0;
  assign isNaNOut = T309 | notSigNaN_invalid;
  assign T309 = T310 | isNaNC;
  assign T310 = isNaNA | isNaNB;
  assign T311 = T312 | isNaNOut;
  assign T312 = totalUnderflowY & roundMagUp;
  assign totalUnderflowY = T317 & T313;
  assign T313 = T316 | T314;
  assign T314 = T315 < 9'h6b;
  assign T315 = sExpY[4'h8:1'h0];
  assign T316 = sExpY[4'h9];
  assign T317 = isZeroY ^ 1'h1;
  assign expOut = T319 | T318;
  assign T318 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T319 = T324 | T320;
  assign T320 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = T322 | T321;
  assign T321 = overflow & overflowY_roundMagUp;
  assign T322 = T323 | isInfC;
  assign T323 = isInfA | isInfB;
  assign T324 = T326 | T325;
  assign T325 = pegMaxFiniteMagOut ? 9'h17f : 9'h0;
  assign T326 = T329 | T327;
  assign T327 = pegMinFiniteMagOut ? 9'h6b : 9'h0;
  assign pegMinFiniteMagOut = T328 & roundMagUp;
  assign T328 = commonCase & totalUnderflowY;
  assign T329 = T332 & T330;
  assign T330 = ~ T331;
  assign T331 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T332 = T335 & T333;
  assign T333 = ~ T334;
  assign T334 = pegMaxFiniteMagOut ? 9'h80 : 9'h0;
  assign T335 = T338 & T336;
  assign T336 = ~ T337;
  assign T337 = pegMinFiniteMagOut ? 9'h194 : 9'h0;
  assign T338 = expY & T339;
  assign T339 = ~ T340;
  assign T340 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign notSpecial_isZeroOut = T341 | totalUnderflowY;
  assign T341 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'h8:1'h0];
  assign signOut = T343 | T342;
  assign T342 = commonCase & signY;
  assign T343 = T358 & uncommonCaseSignOut;
  assign uncommonCaseSignOut = T348 | T344;
  assign T344 = T345 & roundingMode_min;
  assign T345 = T346 & doSubMags;
  assign T346 = T347 & notSpecial_addZeros;
  assign T347 = mulSpecial ^ 1'h1;
  assign T348 = T352 | T349;
  assign T349 = T350 & io_fromPreMul_opSignC;
  assign T350 = T351 & isSpecialC;
  assign T351 = mulSpecial ^ 1'h1;
  assign T352 = T356 | T353;
  assign T353 = T354 & io_fromPreMul_signProd;
  assign T354 = mulSpecial & T355;
  assign T355 = isSpecialC ^ 1'h1;
  assign T356 = T357 & io_fromPreMul_opSignC;
  assign T357 = doSubMags ^ 1'h1;
  assign T358 = isNaNOut ^ 1'h1;
endmodule

module MulAddRecFN_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[48:0] T0;
  wire[48:0] T1;
  wire[48:0] T3;
  wire[47:0] T2;
  wire[23:0] mulAddRecFN_preMul_io_mulAddA;
  wire[23:0] mulAddRecFN_preMul_io_mulAddB;
  wire[47:0] mulAddRecFN_preMul_io_mulAddC;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire mulAddRecFN_preMul_io_toPostMul_signProd;
  wire mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire[6:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire[25:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire[10:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire[1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire[32:0] mulAddRecFN_postMul_io_out;
  wire[4:0] mulAddRecFN_postMul_io_exceptionFlags;


  assign T0 = T3 + T1;
  assign T1 = {1'h0, mulAddRecFN_preMul_io_mulAddC};
  assign T3 = {1'h0, T2};
  assign T2 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign io_out = mulAddRecFN_postMul_io_out;
  MulAddRecFN_preMul_0 mulAddRecFN_preMul(
       .io_op( io_op ),
       .io_a( io_a ),
       .io_b( io_b ),
       .io_c( io_c ),
       .io_roundingMode( io_roundingMode ),
       .io_mulAddA( mulAddRecFN_preMul_io_mulAddA ),
       .io_mulAddB( mulAddRecFN_preMul_io_mulAddB ),
       .io_mulAddC( mulAddRecFN_preMul_io_mulAddC ),
       .io_toPostMul_highExpA( mulAddRecFN_preMul_io_toPostMul_highExpA ),
       .io_toPostMul_isNaN_isQuietNaNA( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA ),
       .io_toPostMul_highExpB( mulAddRecFN_preMul_io_toPostMul_highExpB ),
       .io_toPostMul_isNaN_isQuietNaNB( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB ),
       .io_toPostMul_signProd( mulAddRecFN_preMul_io_toPostMul_signProd ),
       .io_toPostMul_isZeroProd( mulAddRecFN_preMul_io_toPostMul_isZeroProd ),
       .io_toPostMul_opSignC( mulAddRecFN_preMul_io_toPostMul_opSignC ),
       .io_toPostMul_highExpC( mulAddRecFN_preMul_io_toPostMul_highExpC ),
       .io_toPostMul_isNaN_isQuietNaNC( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC ),
       .io_toPostMul_isCDominant( mulAddRecFN_preMul_io_toPostMul_isCDominant ),
       .io_toPostMul_CAlignDist_0( mulAddRecFN_preMul_io_toPostMul_CAlignDist_0 ),
       .io_toPostMul_CAlignDist( mulAddRecFN_preMul_io_toPostMul_CAlignDist ),
       .io_toPostMul_bit0AlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC ),
       .io_toPostMul_highAlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC ),
       .io_toPostMul_sExpSum( mulAddRecFN_preMul_io_toPostMul_sExpSum ),
       .io_toPostMul_roundingMode( mulAddRecFN_preMul_io_toPostMul_roundingMode )
  );
  MulAddRecFN_postMul_0 mulAddRecFN_postMul(
       .io_fromPreMul_highExpA( mulAddRecFN_preMul_io_toPostMul_highExpA ),
       .io_fromPreMul_isNaN_isQuietNaNA( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA ),
       .io_fromPreMul_highExpB( mulAddRecFN_preMul_io_toPostMul_highExpB ),
       .io_fromPreMul_isNaN_isQuietNaNB( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB ),
       .io_fromPreMul_signProd( mulAddRecFN_preMul_io_toPostMul_signProd ),
       .io_fromPreMul_isZeroProd( mulAddRecFN_preMul_io_toPostMul_isZeroProd ),
       .io_fromPreMul_opSignC( mulAddRecFN_preMul_io_toPostMul_opSignC ),
       .io_fromPreMul_highExpC( mulAddRecFN_preMul_io_toPostMul_highExpC ),
       .io_fromPreMul_isNaN_isQuietNaNC( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC ),
       .io_fromPreMul_isCDominant( mulAddRecFN_preMul_io_toPostMul_isCDominant ),
       .io_fromPreMul_CAlignDist_0( mulAddRecFN_preMul_io_toPostMul_CAlignDist_0 ),
       .io_fromPreMul_CAlignDist( mulAddRecFN_preMul_io_toPostMul_CAlignDist ),
       .io_fromPreMul_bit0AlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC ),
       .io_fromPreMul_highAlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC ),
       .io_fromPreMul_sExpSum( mulAddRecFN_preMul_io_toPostMul_sExpSum ),
       .io_fromPreMul_roundingMode( mulAddRecFN_preMul_io_toPostMul_roundingMode ),
       .io_mulAddResult( T0 ),
       .io_out( mulAddRecFN_postMul_io_out ),
       .io_exceptionFlags( mulAddRecFN_postMul_io_exceptionFlags )
  );
endmodule

module FPUFMAPipe_0(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap12,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_div,
    input  io_in_bits_sqrt,
    input  io_in_bits_round,
    input  io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T26;
  reg [2:0] in_rm;
  wire[2:0] T0;
  wire[32:0] T27;
  reg [64:0] in_in3;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[64:0] T28;
  wire[32:0] zero;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[32:0] T29;
  reg [64:0] in_in2;
  wire[64:0] T9;
  wire[64:0] T10;
  wire T11;
  wire[32:0] T30;
  reg [64:0] in_in1;
  wire[64:0] T12;
  wire[1:0] T31;
  reg [4:0] in_cmd;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T32;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [4:0] R20;
  wire[4:0] T21;
  wire[4:0] res_exc;
  reg  valid;
  reg [64:0] R22;
  wire[64:0] T23;
  wire[64:0] res_data;
  wire[64:0] T24;
  reg  R25;
  wire T33;
  wire[32:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R20 = {1{$random}};
    valid = {1{$random}};
    R22 = {3{$random}};
    R25 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T26 = in_rm[1'h1:1'h0];
  assign T0 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T27 = in_in3[6'h20:1'h0];
  assign T1 = T6 ? T28 : T2;
  assign T2 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T28 = {32'h0, zero};
  assign zero = T3 << 6'h20;
  assign T3 = T5 ^ T4;
  assign T4 = io_in_bits_in2[6'h20];
  assign T5 = io_in_bits_in1[6'h20];
  assign T6 = io_in_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T29 = in_in2[6'h20:1'h0];
  assign T9 = T11 ? 65'h80000000 : T10;
  assign T10 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T11 = io_in_valid & io_in_bits_swap23;
  assign T30 = in_in1[6'h20:1'h0];
  assign T12 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T31 = in_cmd[1'h1:1'h0];
  assign T13 = io_in_valid ? T32 : T14;
  assign T14 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T32 = {3'h0, T15};
  assign T15 = {T17, T16};
  assign T16 = io_in_bits_cmd[1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = io_in_bits_cmd[1'h1];
  assign io_out_bits_exc = R20;
  assign T21 = valid ? res_exc : R20;
  assign res_exc = fma_io_exceptionFlags;
  assign io_out_bits_data = R22;
  assign T23 = valid ? res_data : R22;
  assign res_data = T24;
  assign T24 = {32'hffffffff, fma_io_out};
  assign io_out_valid = R25;
  assign T33 = reset ? 1'h0 : valid;
  MulAddRecFN_0 fma(
       .io_op( T31 ),
       .io_a( T30 ),
       .io_b( T29 ),
       .io_c( T27 ),
       .io_roundingMode( T26 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T6) begin
      in_in3 <= T28;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T11) begin
      in_in2 <= 65'h80000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T32;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(valid) begin
      R20 <= res_exc;
    end
    valid <= io_in_valid;
    if(valid) begin
      R22 <= res_data;
    end
    if(reset) begin
      R25 <= 1'h0;
    end else begin
      R25 <= valid;
    end
  end
endmodule

module MulAddRecFN_preMul_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[52:0] io_mulAddA,
    output[52:0] io_mulAddB,
    output[105:0] io_mulAddC,
    output[2:0] io_toPostMul_highExpA,
    output io_toPostMul_isNaN_isQuietNaNA,
    output[2:0] io_toPostMul_highExpB,
    output io_toPostMul_isNaN_isQuietNaNB,
    output io_toPostMul_signProd,
    output io_toPostMul_isZeroProd,
    output io_toPostMul_opSignC,
    output[2:0] io_toPostMul_highExpC,
    output io_toPostMul_isNaN_isQuietNaNC,
    output io_toPostMul_isCDominant,
    output io_toPostMul_CAlignDist_0,
    output[7:0] io_toPostMul_CAlignDist,
    output io_toPostMul_bit0AlignedNegSigC,
    output[54:0] io_toPostMul_highAlignedNegSigC,
    output[13:0] io_toPostMul_sExpSum,
    output[1:0] io_toPostMul_roundingMode
);

  wire[13:0] sExpSum;
  wire[13:0] sExpAlignedProd;
  wire[13:0] T0;
  wire[13:0] T1;
  wire[10:0] T2;
  wire[11:0] expB;
  wire[2:0] T3;
  wire[2:0] T119;
  wire T4;
  wire T5;
  wire[13:0] T120;
  wire[11:0] expA;
  wire[13:0] T121;
  wire[11:0] expC;
  wire CAlignDist_floor;
  wire T6;
  wire[13:0] sNatCAlignDist;
  wire[13:0] T122;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T7;
  wire isZeroA;
  wire[2:0] T8;
  wire[54:0] T9;
  wire[161:0] alignedNegSigC;
  wire[162:0] T10;
  wire T11;
  wire doSubMags;
  wire opSignC;
  wire T12;
  wire T13;
  wire signProd;
  wire T14;
  wire T15;
  wire signB;
  wire signA;
  wire T16;
  wire[52:0] T17;
  wire[52:0] CExtraMask;
  wire[20:0] T18;
  wire[4:0] T19;
  wire T20;
  wire[4:0] T21;
  wire[20:0] T22;
  wire[52:0] T23;
  wire[256:0] T24;
  wire[7:0] CAlignDist;
  wire[7:0] T25;
  wire[7:0] T26;
  wire T27;
  wire[12:0] T28;
  wire[3:0] T29;
  wire[1:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[3:0] T33;
  wire T34;
  wire[1:0] T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire[15:0] T39;
  wire[15:0] T40;
  wire[15:0] T41;
  wire[14:0] T42;
  wire[15:0] T43;
  wire[15:0] T44;
  wire[15:0] T45;
  wire[13:0] T46;
  wire[15:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[11:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[7:0] T54;
  wire[15:0] T55;
  wire[15:0] T56;
  wire[15:0] T123;
  wire[7:0] T57;
  wire[15:0] T58;
  wire[15:0] T124;
  wire[11:0] T59;
  wire[15:0] T60;
  wire[15:0] T125;
  wire[13:0] T61;
  wire[15:0] T62;
  wire[15:0] T126;
  wire[14:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[31:0] T66;
  wire[30:0] T67;
  wire[31:0] T68;
  wire[31:0] T69;
  wire[31:0] T70;
  wire[29:0] T71;
  wire[31:0] T72;
  wire[31:0] T73;
  wire[31:0] T74;
  wire[27:0] T75;
  wire[31:0] T76;
  wire[31:0] T77;
  wire[31:0] T78;
  wire[23:0] T79;
  wire[31:0] T80;
  wire[31:0] T81;
  wire[31:0] T82;
  wire[15:0] T83;
  wire[31:0] T84;
  wire[31:0] T85;
  wire[31:0] T127;
  wire[15:0] T86;
  wire[31:0] T87;
  wire[31:0] T128;
  wire[23:0] T88;
  wire[31:0] T89;
  wire[31:0] T129;
  wire[27:0] T90;
  wire[31:0] T91;
  wire[31:0] T130;
  wire[29:0] T92;
  wire[31:0] T93;
  wire[31:0] T131;
  wire[30:0] T94;
  wire[52:0] sigC;
  wire[51:0] fractC;
  wire T95;
  wire isZeroC;
  wire[2:0] T96;
  wire[161:0] T97;
  wire[161:0] T98;
  wire[161:0] T99;
  wire[160:0] T100;
  wire[107:0] T101;
  wire[107:0] T132;
  wire[52:0] negSigC;
  wire[52:0] T102;
  wire T103;
  wire CAlignDist_0;
  wire T104;
  wire[12:0] T105;
  wire isCDominant;
  wire T106;
  wire T107;
  wire[12:0] T108;
  wire T109;
  wire T110;
  wire[2:0] T111;
  wire T112;
  wire[51:0] fractB;
  wire[2:0] T113;
  wire T114;
  wire[51:0] fractA;
  wire[2:0] T115;
  wire[105:0] T116;
  wire[52:0] sigB;
  wire T117;
  wire[52:0] sigA;
  wire T118;


  assign io_toPostMul_roundingMode = io_roundingMode;
  assign io_toPostMul_sExpSum = sExpSum;
  assign sExpSum = CAlignDist_floor ? T121 : sExpAlignedProd;
  assign sExpAlignedProd = T0 + 14'h38;
  assign T0 = T120 + T1;
  assign T1 = {T3, T2};
  assign T2 = expB[4'ha:1'h0];
  assign expB = io_b[6'h3f:6'h34];
  assign T3 = 3'h0 - T119;
  assign T119 = {2'h0, T4};
  assign T4 = T5 ^ 1'h1;
  assign T5 = expB[4'hb];
  assign T120 = {2'h0, expA};
  assign expA = io_a[6'h3f:6'h34];
  assign T121 = {2'h0, expC};
  assign expC = io_c[6'h3f:6'h34];
  assign CAlignDist_floor = isZeroProd | T6;
  assign T6 = sNatCAlignDist[4'hd];
  assign sNatCAlignDist = sExpAlignedProd - T122;
  assign T122 = {2'h0, expC};
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T7 == 3'h0;
  assign T7 = expB[4'hb:4'h9];
  assign isZeroA = T8 == 3'h0;
  assign T8 = expA[4'hb:4'h9];
  assign io_toPostMul_highAlignedNegSigC = T9;
  assign T9 = alignedNegSigC[8'ha1:7'h6b];
  assign alignedNegSigC = T10[8'ha1:1'h0];
  assign T10 = {T97, T11};
  assign T11 = T16 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T13 ^ T12;
  assign T12 = io_op[1'h0];
  assign T13 = io_c[7'h40];
  assign signProd = T15 ^ T14;
  assign T14 = io_op[1'h1];
  assign T15 = signA ^ signB;
  assign signB = io_b[7'h40];
  assign signA = io_a[7'h40];
  assign T16 = T17 != 53'h0;
  assign T17 = sigC & CExtraMask;
  assign CExtraMask = {T64, T18};
  assign T18 = {T39, T19};
  assign T19 = {T29, T20};
  assign T20 = T21[3'h4];
  assign T21 = T22[5'h14:5'h10];
  assign T22 = T23[6'h34:6'h20];
  assign T23 = T24[8'h93:7'h5f];
  assign T24 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = CAlignDist_floor ? 8'h0 : T25;
  assign T25 = T27 ? T26 : 8'ha1;
  assign T26 = sNatCAlignDist[3'h7:1'h0];
  assign T27 = T28 < 13'ha1;
  assign T28 = sNatCAlignDist[4'hc:1'h0];
  assign T29 = {T35, T30};
  assign T30 = {T34, T31};
  assign T31 = T32[1'h1];
  assign T32 = T33[2'h3:2'h2];
  assign T33 = T21[2'h3:1'h0];
  assign T34 = T32[1'h0];
  assign T35 = {T38, T36};
  assign T36 = T37[1'h1];
  assign T37 = T33[1'h1:1'h0];
  assign T38 = T37[1'h0];
  assign T39 = T62 | T40;
  assign T40 = T41 & 16'haaaa;
  assign T41 = T42 << 1'h1;
  assign T42 = T43[4'he:1'h0];
  assign T43 = T60 | T44;
  assign T44 = T45 & 16'hcccc;
  assign T45 = T46 << 2'h2;
  assign T46 = T47[4'hd:1'h0];
  assign T47 = T58 | T48;
  assign T48 = T49 & 16'hf0f0;
  assign T49 = T50 << 3'h4;
  assign T50 = T51[4'hb:1'h0];
  assign T51 = T56 | T52;
  assign T52 = T53 & 16'hff00;
  assign T53 = T54 << 4'h8;
  assign T54 = T55[3'h7:1'h0];
  assign T55 = T22[4'hf:1'h0];
  assign T56 = T123 & 16'hff;
  assign T123 = {8'h0, T57};
  assign T57 = T55 >> 4'h8;
  assign T58 = T124 & 16'hf0f;
  assign T124 = {4'h0, T59};
  assign T59 = T51 >> 3'h4;
  assign T60 = T125 & 16'h3333;
  assign T125 = {2'h0, T61};
  assign T61 = T47 >> 2'h2;
  assign T62 = T126 & 16'h5555;
  assign T126 = {1'h0, T63};
  assign T63 = T43 >> 1'h1;
  assign T64 = T93 | T65;
  assign T65 = T66 & 32'haaaaaaaa;
  assign T66 = T67 << 1'h1;
  assign T67 = T68[5'h1e:1'h0];
  assign T68 = T91 | T69;
  assign T69 = T70 & 32'hcccccccc;
  assign T70 = T71 << 2'h2;
  assign T71 = T72[5'h1d:1'h0];
  assign T72 = T89 | T73;
  assign T73 = T74 & 32'hf0f0f0f0;
  assign T74 = T75 << 3'h4;
  assign T75 = T76[5'h1b:1'h0];
  assign T76 = T87 | T77;
  assign T77 = T78 & 32'hff00ff00;
  assign T78 = T79 << 4'h8;
  assign T79 = T80[5'h17:1'h0];
  assign T80 = T85 | T81;
  assign T81 = T82 & 32'hffff0000;
  assign T82 = T83 << 5'h10;
  assign T83 = T84[4'hf:1'h0];
  assign T84 = T23[5'h1f:1'h0];
  assign T85 = T127 & 32'hffff;
  assign T127 = {16'h0, T86};
  assign T86 = T84 >> 5'h10;
  assign T87 = T128 & 32'hff00ff;
  assign T128 = {8'h0, T88};
  assign T88 = T80 >> 4'h8;
  assign T89 = T129 & 32'hf0f0f0f;
  assign T129 = {4'h0, T90};
  assign T90 = T76 >> 3'h4;
  assign T91 = T130 & 32'h33333333;
  assign T130 = {2'h0, T92};
  assign T92 = T72 >> 2'h2;
  assign T93 = T131 & 32'h55555555;
  assign T131 = {1'h0, T94};
  assign T94 = T68 >> 1'h1;
  assign sigC = {T95, fractC};
  assign fractC = io_c[6'h33:1'h0];
  assign T95 = isZeroC ^ 1'h1;
  assign isZeroC = T96 == 3'h0;
  assign T96 = expC[4'hb:4'h9];
  assign T97 = $signed(T98) >>> CAlignDist;
  assign T98 = T99;
  assign T99 = {doSubMags, T100};
  assign T100 = {negSigC, T101};
  assign T101 = 108'h0 - T132;
  assign T132 = {107'h0, doSubMags};
  assign negSigC = doSubMags ? T102 : sigC;
  assign T102 = ~ sigC;
  assign io_toPostMul_bit0AlignedNegSigC = T103;
  assign T103 = alignedNegSigC[1'h0];
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign CAlignDist_0 = CAlignDist_floor | T104;
  assign T104 = T105 == 13'h0;
  assign T105 = sNatCAlignDist[4'hc:1'h0];
  assign io_toPostMul_isCDominant = isCDominant;
  assign isCDominant = T109 & T106;
  assign T106 = CAlignDist_floor | T107;
  assign T107 = T108 < 13'h36;
  assign T108 = sNatCAlignDist[4'hc:1'h0];
  assign T109 = isZeroC ^ 1'h1;
  assign io_toPostMul_isNaN_isQuietNaNC = T110;
  assign T110 = fractC[6'h33];
  assign io_toPostMul_highExpC = T111;
  assign T111 = expC[4'hb:4'h9];
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isNaN_isQuietNaNB = T112;
  assign T112 = fractB[6'h33];
  assign fractB = io_b[6'h33:1'h0];
  assign io_toPostMul_highExpB = T113;
  assign T113 = expB[4'hb:4'h9];
  assign io_toPostMul_isNaN_isQuietNaNA = T114;
  assign T114 = fractA[6'h33];
  assign fractA = io_a[6'h33:1'h0];
  assign io_toPostMul_highExpA = T115;
  assign T115 = expA[4'hb:4'h9];
  assign io_mulAddC = T116;
  assign T116 = alignedNegSigC[7'h6a:1'h1];
  assign io_mulAddB = sigB;
  assign sigB = {T117, fractB};
  assign T117 = isZeroB ^ 1'h1;
  assign io_mulAddA = sigA;
  assign sigA = {T118, fractA};
  assign T118 = isZeroA ^ 1'h1;
endmodule

module MulAddRecFN_postMul_1(
    input [2:0] io_fromPreMul_highExpA,
    input  io_fromPreMul_isNaN_isQuietNaNA,
    input [2:0] io_fromPreMul_highExpB,
    input  io_fromPreMul_isNaN_isQuietNaNB,
    input  io_fromPreMul_signProd,
    input  io_fromPreMul_isZeroProd,
    input  io_fromPreMul_opSignC,
    input [2:0] io_fromPreMul_highExpC,
    input  io_fromPreMul_isNaN_isQuietNaNC,
    input  io_fromPreMul_isCDominant,
    input  io_fromPreMul_CAlignDist_0,
    input [7:0] io_fromPreMul_CAlignDist,
    input  io_fromPreMul_bit0AlignedNegSigC,
    input [54:0] io_fromPreMul_highAlignedNegSigC,
    input [13:0] io_fromPreMul_sExpSum,
    input [1:0] io_fromPreMul_roundingMode,
    input [106:0] io_mulAddResult,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[56:0] T4;
  wire[56:0] T431;
  wire[54:0] T5;
  wire[55:0] roundMask;
  wire[55:0] T6;
  wire[53:0] T7;
  wire[53:0] T432;
  wire T8;
  wire[53:0] T9;
  wire[21:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[5:0] T15;
  wire[21:0] T16;
  wire[53:0] T17;
  wire[8192:0] T18;
  wire[12:0] T19;
  wire[12:0] sExpX3_13;
  wire[13:0] sExpX3;
  wire[13:0] T433;
  wire[7:0] estNormDist;
  wire[7:0] T20;
  wire[7:0] estNormNeg_dist;
  wire[7:0] T434;
  wire[6:0] T435;
  wire[6:0] T436;
  wire[6:0] T437;
  wire[6:0] T438;
  wire[6:0] T439;
  wire[6:0] T440;
  wire[6:0] T441;
  wire[6:0] T442;
  wire[6:0] T443;
  wire[6:0] T444;
  wire[6:0] T445;
  wire[6:0] T446;
  wire[6:0] T447;
  wire[6:0] T448;
  wire[6:0] T449;
  wire[6:0] T450;
  wire[6:0] T451;
  wire[6:0] T452;
  wire[6:0] T453;
  wire[6:0] T454;
  wire[6:0] T455;
  wire[6:0] T456;
  wire[6:0] T457;
  wire[6:0] T458;
  wire[6:0] T459;
  wire[6:0] T460;
  wire[6:0] T461;
  wire[6:0] T462;
  wire[6:0] T463;
  wire[6:0] T464;
  wire[6:0] T465;
  wire[6:0] T466;
  wire[6:0] T467;
  wire[6:0] T468;
  wire[6:0] T469;
  wire[6:0] T470;
  wire[6:0] T471;
  wire[6:0] T472;
  wire[6:0] T473;
  wire[6:0] T474;
  wire[6:0] T475;
  wire[6:0] T476;
  wire[6:0] T477;
  wire[6:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[5:0] T493;
  wire[5:0] T494;
  wire[5:0] T495;
  wire[5:0] T496;
  wire[5:0] T497;
  wire[5:0] T498;
  wire[5:0] T499;
  wire[5:0] T500;
  wire[5:0] T501;
  wire[5:0] T502;
  wire[5:0] T503;
  wire[5:0] T504;
  wire[5:0] T505;
  wire[5:0] T506;
  wire[5:0] T507;
  wire[5:0] T508;
  wire[5:0] T509;
  wire[5:0] T510;
  wire[4:0] T511;
  wire[4:0] T512;
  wire[4:0] T513;
  wire[4:0] T514;
  wire[4:0] T515;
  wire[4:0] T516;
  wire[4:0] T517;
  wire[4:0] T518;
  wire[4:0] T519;
  wire[4:0] T520;
  wire[4:0] T521;
  wire[4:0] T522;
  wire[4:0] T523;
  wire[4:0] T524;
  wire[4:0] T525;
  wire[4:0] T526;
  wire[3:0] T527;
  wire[3:0] T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[3:0] T532;
  wire[3:0] T533;
  wire[3:0] T534;
  wire[2:0] T535;
  wire[2:0] T536;
  wire[2:0] T537;
  wire[2:0] T538;
  wire[1:0] T539;
  wire[1:0] T540;
  wire T541;
  wire[107:0] T22;
  wire[107:0] T23;
  wire[108:0] T24;
  wire[108:0] T25;
  wire[107:0] T26;
  wire[107:0] T27;
  wire[161:0] sigSum;
  wire[106:0] T28;
  wire[105:0] T29;
  wire[54:0] T30;
  wire[54:0] T31;
  wire T32;
  wire[108:0] T542;
  wire[107:0] T33;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire notCDom_signSigSum;
  wire[7:0] CDom_estNormDist;
  wire[7:0] T649;
  wire[5:0] T34;
  wire[7:0] T35;
  wire T36;
  wire doSubMags;
  wire T37;
  wire[3:0] T38;
  wire[1:0] T39;
  wire T40;
  wire[1:0] T41;
  wire[3:0] T42;
  wire T43;
  wire[1:0] T44;
  wire T45;
  wire[1:0] T46;
  wire T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[15:0] T50;
  wire[14:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[15:0] T54;
  wire[13:0] T55;
  wire[15:0] T56;
  wire[15:0] T57;
  wire[15:0] T58;
  wire[11:0] T59;
  wire[15:0] T60;
  wire[15:0] T61;
  wire[15:0] T62;
  wire[7:0] T63;
  wire[15:0] T64;
  wire[15:0] T65;
  wire[15:0] T650;
  wire[7:0] T66;
  wire[15:0] T67;
  wire[15:0] T651;
  wire[11:0] T68;
  wire[15:0] T69;
  wire[15:0] T652;
  wire[13:0] T70;
  wire[15:0] T71;
  wire[15:0] T653;
  wire[14:0] T72;
  wire[31:0] T73;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[30:0] T76;
  wire[31:0] T77;
  wire[31:0] T78;
  wire[31:0] T79;
  wire[29:0] T80;
  wire[31:0] T81;
  wire[31:0] T82;
  wire[31:0] T83;
  wire[27:0] T84;
  wire[31:0] T85;
  wire[31:0] T86;
  wire[31:0] T87;
  wire[23:0] T88;
  wire[31:0] T89;
  wire[31:0] T90;
  wire[31:0] T91;
  wire[15:0] T92;
  wire[31:0] T93;
  wire[31:0] T94;
  wire[31:0] T654;
  wire[15:0] T95;
  wire[31:0] T96;
  wire[31:0] T655;
  wire[23:0] T97;
  wire[31:0] T98;
  wire[31:0] T656;
  wire[27:0] T99;
  wire[31:0] T100;
  wire[31:0] T657;
  wire[29:0] T101;
  wire[31:0] T102;
  wire[31:0] T658;
  wire[30:0] T103;
  wire[55:0] T104;
  wire[55:0] T659;
  wire T105;
  wire[56:0] sigX3;
  wire[87:0] T106;
  wire T107;
  wire T108;
  wire[31:0] T109;
  wire[31:0] absSigSumExtraMask;
  wire[30:0] T110;
  wire[14:0] T111;
  wire[6:0] T112;
  wire[2:0] T113;
  wire T114;
  wire[2:0] T115;
  wire[6:0] T116;
  wire[14:0] T117;
  wire[30:0] T118;
  wire[32:0] T119;
  wire[4:0] normTo2ShiftDist;
  wire[4:0] estNormDist_5;
  wire[1:0] T120;
  wire T121;
  wire[1:0] T122;
  wire T123;
  wire[3:0] T124;
  wire[1:0] T125;
  wire T126;
  wire[1:0] T127;
  wire[3:0] T128;
  wire T129;
  wire[1:0] T130;
  wire T131;
  wire[1:0] T132;
  wire T133;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[6:0] T137;
  wire[7:0] T138;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[5:0] T141;
  wire[7:0] T142;
  wire[7:0] T143;
  wire[7:0] T144;
  wire[3:0] T145;
  wire[7:0] T146;
  wire[7:0] T147;
  wire[7:0] T660;
  wire[3:0] T148;
  wire[7:0] T149;
  wire[7:0] T661;
  wire[5:0] T150;
  wire[7:0] T151;
  wire[7:0] T662;
  wire[6:0] T152;
  wire[15:0] T153;
  wire[15:0] T154;
  wire[15:0] T155;
  wire[14:0] T156;
  wire[15:0] T157;
  wire[15:0] T158;
  wire[15:0] T159;
  wire[13:0] T160;
  wire[15:0] T161;
  wire[15:0] T162;
  wire[15:0] T163;
  wire[11:0] T164;
  wire[15:0] T165;
  wire[15:0] T166;
  wire[15:0] T167;
  wire[7:0] T168;
  wire[15:0] T169;
  wire[15:0] T170;
  wire[15:0] T663;
  wire[7:0] T171;
  wire[15:0] T172;
  wire[15:0] T664;
  wire[11:0] T173;
  wire[15:0] T174;
  wire[15:0] T665;
  wire[13:0] T175;
  wire[15:0] T176;
  wire[15:0] T666;
  wire[14:0] T177;
  wire[31:0] T178;
  wire[87:0] cFirstNormAbsSigSum;
  wire[87:0] T667;
  wire[86:0] T179;
  wire[86:0] notCDom_pos_firstNormAbsSigSum;
  wire[86:0] T180;
  wire[86:0] T181;
  wire[53:0] T182;
  wire[53:0] T668;
  wire[32:0] T183;
  wire[86:0] T184;
  wire[86:0] T185;
  wire[85:0] T186;
  wire[85:0] T669;
  wire T187;
  wire[86:0] T670;
  wire[65:0] T188;
  wire T189;
  wire T190;
  wire[1:0] firstReduceSigSum;
  wire T191;
  wire[43:0] T192;
  wire T193;
  wire[31:0] T194;
  wire T195;
  wire T196;
  wire[1:0] firstReduceComplSigSum;
  wire T197;
  wire[43:0] T198;
  wire[161:0] complSigSum;
  wire T199;
  wire[31:0] T200;
  wire[64:0] T201;
  wire T202;
  wire T203;
  wire[86:0] T204;
  wire[86:0] T205;
  wire T206;
  wire T207;
  wire[10:0] T208;
  wire T209;
  wire[10:0] T210;
  wire[85:0] T211;
  wire[86:0] T212;
  wire[21:0] T213;
  wire[21:0] T671;
  wire[64:0] T214;
  wire T215;
  wire T216;
  wire[86:0] CDom_firstNormAbsSigSum;
  wire[86:0] T217;
  wire[86:0] T218;
  wire T219;
  wire[85:0] T220;
  wire T221;
  wire T222;
  wire[86:0] T223;
  wire[86:0] T224;
  wire[86:0] T225;
  wire T226;
  wire[85:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire[86:0] T231;
  wire[86:0] T232;
  wire[86:0] T233;
  wire T234;
  wire[85:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire[86:0] T239;
  wire[86:0] T240;
  wire T241;
  wire[85:0] T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[87:0] T247;
  wire[87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[87:0] T248;
  wire[87:0] T249;
  wire[33:0] T250;
  wire[87:0] T251;
  wire[87:0] T252;
  wire[1:0] T253;
  wire[87:0] T672;
  wire[64:0] T254;
  wire T255;
  wire[63:0] T256;
  wire T257;
  wire T258;
  wire[87:0] T259;
  wire[87:0] T260;
  wire T261;
  wire[10:0] T262;
  wire[86:0] T263;
  wire[87:0] T264;
  wire[65:0] T265;
  wire T266;
  wire T267;
  wire[87:0] T673;
  wire T268;
  wire[31:0] T269;
  wire[31:0] T270;
  wire[31:0] T271;
  wire[86:0] T272;
  wire[86:0] T273;
  wire roundPosBit;
  wire[56:0] T274;
  wire[56:0] T674;
  wire[55:0] roundPosMask;
  wire[55:0] T675;
  wire[54:0] T275;
  wire[54:0] T276;
  wire T277;
  wire allRound;
  wire allRoundExtra;
  wire[56:0] T278;
  wire[56:0] T676;
  wire[54:0] T279;
  wire[56:0] T280;
  wire doIncrSig;
  wire T281;
  wire T282;
  wire T283;
  wire commonCase;
  wire T284;
  wire notSpecial_addZeros;
  wire isZeroC;
  wire T285;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T286;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T287;
  wire isSpecialA;
  wire[1:0] T288;
  wire underflow;
  wire underflowY;
  wire T289;
  wire T290;
  wire[12:0] T677;
  wire[10:0] T291;
  wire sigX3Shift1;
  wire[1:0] T292;
  wire T293;
  wire overflow;
  wire overflowY;
  wire[2:0] T294;
  wire[13:0] sExpY;
  wire[13:0] T295;
  wire[13:0] T296;
  wire T297;
  wire[1:0] T298;
  wire[54:0] sigY3;
  wire[54:0] T299;
  wire[54:0] T300;
  wire[54:0] T301;
  wire[54:0] T302;
  wire[54:0] roundUp_sigY3;
  wire[54:0] T303;
  wire[54:0] T304;
  wire[56:0] T305;
  wire[56:0] T678;
  wire roundEven;
  wire T306;
  wire T307;
  wire T308;
  wire roundingMode_nearest_even;
  wire T309;
  wire T310;
  wire T311;
  wire[54:0] T312;
  wire[54:0] T313;
  wire roundUp;
  wire T314;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T315;
  wire doNegSignSum;
  wire T316;
  wire T317;
  wire isZeroY;
  wire[2:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[54:0] T332;
  wire[54:0] T333;
  wire[56:0] T334;
  wire[56:0] T679;
  wire[55:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[13:0] T339;
  wire[13:0] T340;
  wire T341;
  wire[13:0] T342;
  wire[13:0] T343;
  wire T344;
  wire[1:0] T345;
  wire invalid;
  wire notSigNaN_invalid;
  wire T346;
  wire T347;
  wire isInfC;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire isInfB;
  wire T352;
  wire T353;
  wire isInfA;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire isNaNB;
  wire T358;
  wire T359;
  wire isNaNA;
  wire T360;
  wire T361;
  wire T362;
  wire isZeroA;
  wire T363;
  wire isZeroB;
  wire T364;
  wire isSigNaNC;
  wire T365;
  wire isNaNC;
  wire T366;
  wire T367;
  wire isSigNaNB;
  wire T368;
  wire isSigNaNA;
  wire T369;
  wire[64:0] T370;
  wire[63:0] T371;
  wire[51:0] fractOut;
  wire[51:0] T372;
  wire[51:0] T680;
  wire pegMaxFiniteMagOut;
  wire T373;
  wire overflowY_roundMagUp;
  wire roundMagUp;
  wire T374;
  wire T375;
  wire T376;
  wire[51:0] T377;
  wire[51:0] fractY;
  wire[51:0] T378;
  wire[51:0] T379;
  wire[51:0] T380;
  wire isNaNOut;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire totalUnderflowY;
  wire T385;
  wire T386;
  wire[11:0] T387;
  wire T388;
  wire T389;
  wire[11:0] expOut;
  wire[11:0] T390;
  wire[11:0] T391;
  wire[11:0] T392;
  wire notNaN_isInfOut;
  wire T393;
  wire T394;
  wire T395;
  wire[11:0] T396;
  wire[11:0] T397;
  wire[11:0] T398;
  wire[11:0] T399;
  wire pegMinFiniteMagOut;
  wire T400;
  wire[11:0] T401;
  wire[11:0] T402;
  wire[11:0] T403;
  wire[11:0] T404;
  wire[11:0] T405;
  wire[11:0] T406;
  wire[11:0] T407;
  wire[11:0] T408;
  wire[11:0] T409;
  wire[11:0] T410;
  wire[11:0] T411;
  wire[11:0] T412;
  wire notSpecial_isZeroOut;
  wire T413;
  wire[11:0] expY;
  wire signOut;
  wire T414;
  wire T415;
  wire uncommonCaseSignOut;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;


  assign io_exceptionFlags = T0;
  assign T0 = {T345, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T277 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 57'h0;
  assign T4 = sigX3 & T431;
  assign T431 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T104 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T432;
  assign T432 = {53'h0, T8};
  assign T8 = sigX3[6'h37];
  assign T9 = {T73, T10};
  assign T10 = {T48, T11};
  assign T11 = {T38, T12};
  assign T12 = {T37, T13};
  assign T13 = T14[1'h1];
  assign T14 = T15[3'h5:3'h4];
  assign T15 = T16[5'h15:5'h10];
  assign T16 = T17[6'h35:6'h20];
  assign T17 = T18[11'h403:10'h3ce];
  assign T18 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T19;
  assign T19 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'hc:1'h0];
  assign sExpX3 = io_fromPreMul_sExpSum - T433;
  assign T433 = {6'h0, estNormDist};
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : T20;
  assign T20 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = 8'ha0 - T434;
  assign T434 = {1'h0, T435};
  assign T435 = T648 ? 7'h6b : T436;
  assign T436 = T647 ? 7'h6a : T437;
  assign T437 = T646 ? 7'h69 : T438;
  assign T438 = T645 ? 7'h68 : T439;
  assign T439 = T644 ? 7'h67 : T440;
  assign T440 = T643 ? 7'h66 : T441;
  assign T441 = T642 ? 7'h65 : T442;
  assign T442 = T641 ? 7'h64 : T443;
  assign T443 = T640 ? 7'h63 : T444;
  assign T444 = T639 ? 7'h62 : T445;
  assign T445 = T638 ? 7'h61 : T446;
  assign T446 = T637 ? 7'h60 : T447;
  assign T447 = T636 ? 7'h5f : T448;
  assign T448 = T635 ? 7'h5e : T449;
  assign T449 = T634 ? 7'h5d : T450;
  assign T450 = T633 ? 7'h5c : T451;
  assign T451 = T632 ? 7'h5b : T452;
  assign T452 = T631 ? 7'h5a : T453;
  assign T453 = T630 ? 7'h59 : T454;
  assign T454 = T629 ? 7'h58 : T455;
  assign T455 = T628 ? 7'h57 : T456;
  assign T456 = T627 ? 7'h56 : T457;
  assign T457 = T626 ? 7'h55 : T458;
  assign T458 = T625 ? 7'h54 : T459;
  assign T459 = T624 ? 7'h53 : T460;
  assign T460 = T623 ? 7'h52 : T461;
  assign T461 = T622 ? 7'h51 : T462;
  assign T462 = T621 ? 7'h50 : T463;
  assign T463 = T620 ? 7'h4f : T464;
  assign T464 = T619 ? 7'h4e : T465;
  assign T465 = T618 ? 7'h4d : T466;
  assign T466 = T617 ? 7'h4c : T467;
  assign T467 = T616 ? 7'h4b : T468;
  assign T468 = T615 ? 7'h4a : T469;
  assign T469 = T614 ? 7'h49 : T470;
  assign T470 = T613 ? 7'h48 : T471;
  assign T471 = T612 ? 7'h47 : T472;
  assign T472 = T611 ? 7'h46 : T473;
  assign T473 = T610 ? 7'h45 : T474;
  assign T474 = T609 ? 7'h44 : T475;
  assign T475 = T608 ? 7'h43 : T476;
  assign T476 = T607 ? 7'h42 : T477;
  assign T477 = T606 ? 7'h41 : T478;
  assign T478 = T605 ? 7'h40 : T479;
  assign T479 = T604 ? 6'h3f : T480;
  assign T480 = T603 ? 6'h3e : T481;
  assign T481 = T602 ? 6'h3d : T482;
  assign T482 = T601 ? 6'h3c : T483;
  assign T483 = T600 ? 6'h3b : T484;
  assign T484 = T599 ? 6'h3a : T485;
  assign T485 = T598 ? 6'h39 : T486;
  assign T486 = T597 ? 6'h38 : T487;
  assign T487 = T596 ? 6'h37 : T488;
  assign T488 = T595 ? 6'h36 : T489;
  assign T489 = T594 ? 6'h35 : T490;
  assign T490 = T593 ? 6'h34 : T491;
  assign T491 = T592 ? 6'h33 : T492;
  assign T492 = T591 ? 6'h32 : T493;
  assign T493 = T590 ? 6'h31 : T494;
  assign T494 = T589 ? 6'h30 : T495;
  assign T495 = T588 ? 6'h2f : T496;
  assign T496 = T587 ? 6'h2e : T497;
  assign T497 = T586 ? 6'h2d : T498;
  assign T498 = T585 ? 6'h2c : T499;
  assign T499 = T584 ? 6'h2b : T500;
  assign T500 = T583 ? 6'h2a : T501;
  assign T501 = T582 ? 6'h29 : T502;
  assign T502 = T581 ? 6'h28 : T503;
  assign T503 = T580 ? 6'h27 : T504;
  assign T504 = T579 ? 6'h26 : T505;
  assign T505 = T578 ? 6'h25 : T506;
  assign T506 = T577 ? 6'h24 : T507;
  assign T507 = T576 ? 6'h23 : T508;
  assign T508 = T575 ? 6'h22 : T509;
  assign T509 = T574 ? 6'h21 : T510;
  assign T510 = T573 ? 6'h20 : T511;
  assign T511 = T572 ? 5'h1f : T512;
  assign T512 = T571 ? 5'h1e : T513;
  assign T513 = T570 ? 5'h1d : T514;
  assign T514 = T569 ? 5'h1c : T515;
  assign T515 = T568 ? 5'h1b : T516;
  assign T516 = T567 ? 5'h1a : T517;
  assign T517 = T566 ? 5'h19 : T518;
  assign T518 = T565 ? 5'h18 : T519;
  assign T519 = T564 ? 5'h17 : T520;
  assign T520 = T563 ? 5'h16 : T521;
  assign T521 = T562 ? 5'h15 : T522;
  assign T522 = T561 ? 5'h14 : T523;
  assign T523 = T560 ? 5'h13 : T524;
  assign T524 = T559 ? 5'h12 : T525;
  assign T525 = T558 ? 5'h11 : T526;
  assign T526 = T557 ? 5'h10 : T527;
  assign T527 = T556 ? 4'hf : T528;
  assign T528 = T555 ? 4'he : T529;
  assign T529 = T554 ? 4'hd : T530;
  assign T530 = T553 ? 4'hc : T531;
  assign T531 = T552 ? 4'hb : T532;
  assign T532 = T551 ? 4'ha : T533;
  assign T533 = T550 ? 4'h9 : T534;
  assign T534 = T549 ? 4'h8 : T535;
  assign T535 = T548 ? 3'h7 : T536;
  assign T536 = T547 ? 3'h6 : T537;
  assign T537 = T546 ? 3'h5 : T538;
  assign T538 = T545 ? 3'h4 : T539;
  assign T539 = T544 ? 2'h3 : T540;
  assign T540 = T543 ? 2'h2 : T541;
  assign T541 = T22[1'h1];
  assign T22 = T23;
  assign T23 = T24[7'h6b:1'h0];
  assign T24 = T542 ^ T25;
  assign T25 = T26 << 1'h1;
  assign T26 = 108'h0 | T27;
  assign T27 = sigSum[7'h6c:1'h1];
  assign sigSum = {T30, T28};
  assign T28 = {T29, io_fromPreMul_bit0AlignedNegSigC};
  assign T29 = io_mulAddResult[7'h69:1'h0];
  assign T30 = T32 ? T31 : io_fromPreMul_highAlignedNegSigC;
  assign T31 = io_fromPreMul_highAlignedNegSigC + 55'h1;
  assign T32 = io_mulAddResult[7'h6a];
  assign T542 = {1'h0, T33};
  assign T33 = 108'h0 ^ T27;
  assign T543 = T22[2'h2];
  assign T544 = T22[2'h3];
  assign T545 = T22[3'h4];
  assign T546 = T22[3'h5];
  assign T547 = T22[3'h6];
  assign T548 = T22[3'h7];
  assign T549 = T22[4'h8];
  assign T550 = T22[4'h9];
  assign T551 = T22[4'ha];
  assign T552 = T22[4'hb];
  assign T553 = T22[4'hc];
  assign T554 = T22[4'hd];
  assign T555 = T22[4'he];
  assign T556 = T22[4'hf];
  assign T557 = T22[5'h10];
  assign T558 = T22[5'h11];
  assign T559 = T22[5'h12];
  assign T560 = T22[5'h13];
  assign T561 = T22[5'h14];
  assign T562 = T22[5'h15];
  assign T563 = T22[5'h16];
  assign T564 = T22[5'h17];
  assign T565 = T22[5'h18];
  assign T566 = T22[5'h19];
  assign T567 = T22[5'h1a];
  assign T568 = T22[5'h1b];
  assign T569 = T22[5'h1c];
  assign T570 = T22[5'h1d];
  assign T571 = T22[5'h1e];
  assign T572 = T22[5'h1f];
  assign T573 = T22[6'h20];
  assign T574 = T22[6'h21];
  assign T575 = T22[6'h22];
  assign T576 = T22[6'h23];
  assign T577 = T22[6'h24];
  assign T578 = T22[6'h25];
  assign T579 = T22[6'h26];
  assign T580 = T22[6'h27];
  assign T581 = T22[6'h28];
  assign T582 = T22[6'h29];
  assign T583 = T22[6'h2a];
  assign T584 = T22[6'h2b];
  assign T585 = T22[6'h2c];
  assign T586 = T22[6'h2d];
  assign T587 = T22[6'h2e];
  assign T588 = T22[6'h2f];
  assign T589 = T22[6'h30];
  assign T590 = T22[6'h31];
  assign T591 = T22[6'h32];
  assign T592 = T22[6'h33];
  assign T593 = T22[6'h34];
  assign T594 = T22[6'h35];
  assign T595 = T22[6'h36];
  assign T596 = T22[6'h37];
  assign T597 = T22[6'h38];
  assign T598 = T22[6'h39];
  assign T599 = T22[6'h3a];
  assign T600 = T22[6'h3b];
  assign T601 = T22[6'h3c];
  assign T602 = T22[6'h3d];
  assign T603 = T22[6'h3e];
  assign T604 = T22[6'h3f];
  assign T605 = T22[7'h40];
  assign T606 = T22[7'h41];
  assign T607 = T22[7'h42];
  assign T608 = T22[7'h43];
  assign T609 = T22[7'h44];
  assign T610 = T22[7'h45];
  assign T611 = T22[7'h46];
  assign T612 = T22[7'h47];
  assign T613 = T22[7'h48];
  assign T614 = T22[7'h49];
  assign T615 = T22[7'h4a];
  assign T616 = T22[7'h4b];
  assign T617 = T22[7'h4c];
  assign T618 = T22[7'h4d];
  assign T619 = T22[7'h4e];
  assign T620 = T22[7'h4f];
  assign T621 = T22[7'h50];
  assign T622 = T22[7'h51];
  assign T623 = T22[7'h52];
  assign T624 = T22[7'h53];
  assign T625 = T22[7'h54];
  assign T626 = T22[7'h55];
  assign T627 = T22[7'h56];
  assign T628 = T22[7'h57];
  assign T629 = T22[7'h58];
  assign T630 = T22[7'h59];
  assign T631 = T22[7'h5a];
  assign T632 = T22[7'h5b];
  assign T633 = T22[7'h5c];
  assign T634 = T22[7'h5d];
  assign T635 = T22[7'h5e];
  assign T636 = T22[7'h5f];
  assign T637 = T22[7'h60];
  assign T638 = T22[7'h61];
  assign T639 = T22[7'h62];
  assign T640 = T22[7'h63];
  assign T641 = T22[7'h64];
  assign T642 = T22[7'h65];
  assign T643 = T22[7'h66];
  assign T644 = T22[7'h67];
  assign T645 = T22[7'h68];
  assign T646 = T22[7'h69];
  assign T647 = T22[7'h6a];
  assign T648 = T22[7'h6b];
  assign notCDom_signSigSum = sigSum[7'h6d];
  assign CDom_estNormDist = T36 ? io_fromPreMul_CAlignDist : T649;
  assign T649 = {2'h0, T34};
  assign T34 = T35[3'h5:1'h0];
  assign T35 = io_fromPreMul_CAlignDist - 8'h1;
  assign T36 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T37 = T14[1'h0];
  assign T38 = {T44, T39};
  assign T39 = {T43, T40};
  assign T40 = T41[1'h1];
  assign T41 = T42[2'h3:2'h2];
  assign T42 = T15[2'h3:1'h0];
  assign T43 = T41[1'h0];
  assign T44 = {T47, T45};
  assign T45 = T46[1'h1];
  assign T46 = T42[1'h1:1'h0];
  assign T47 = T46[1'h0];
  assign T48 = T71 | T49;
  assign T49 = T50 & 16'haaaa;
  assign T50 = T51 << 1'h1;
  assign T51 = T52[4'he:1'h0];
  assign T52 = T69 | T53;
  assign T53 = T54 & 16'hcccc;
  assign T54 = T55 << 2'h2;
  assign T55 = T56[4'hd:1'h0];
  assign T56 = T67 | T57;
  assign T57 = T58 & 16'hf0f0;
  assign T58 = T59 << 3'h4;
  assign T59 = T60[4'hb:1'h0];
  assign T60 = T65 | T61;
  assign T61 = T62 & 16'hff00;
  assign T62 = T63 << 4'h8;
  assign T63 = T64[3'h7:1'h0];
  assign T64 = T16[4'hf:1'h0];
  assign T65 = T650 & 16'hff;
  assign T650 = {8'h0, T66};
  assign T66 = T64 >> 4'h8;
  assign T67 = T651 & 16'hf0f;
  assign T651 = {4'h0, T68};
  assign T68 = T60 >> 3'h4;
  assign T69 = T652 & 16'h3333;
  assign T652 = {2'h0, T70};
  assign T70 = T56 >> 2'h2;
  assign T71 = T653 & 16'h5555;
  assign T653 = {1'h0, T72};
  assign T72 = T52 >> 1'h1;
  assign T73 = T102 | T74;
  assign T74 = T75 & 32'haaaaaaaa;
  assign T75 = T76 << 1'h1;
  assign T76 = T77[5'h1e:1'h0];
  assign T77 = T100 | T78;
  assign T78 = T79 & 32'hcccccccc;
  assign T79 = T80 << 2'h2;
  assign T80 = T81[5'h1d:1'h0];
  assign T81 = T98 | T82;
  assign T82 = T83 & 32'hf0f0f0f0;
  assign T83 = T84 << 3'h4;
  assign T84 = T85[5'h1b:1'h0];
  assign T85 = T96 | T86;
  assign T86 = T87 & 32'hff00ff00;
  assign T87 = T88 << 4'h8;
  assign T88 = T89[5'h17:1'h0];
  assign T89 = T94 | T90;
  assign T90 = T91 & 32'hffff0000;
  assign T91 = T92 << 5'h10;
  assign T92 = T93[4'hf:1'h0];
  assign T93 = T17[5'h1f:1'h0];
  assign T94 = T654 & 32'hffff;
  assign T654 = {16'h0, T95};
  assign T95 = T93 >> 5'h10;
  assign T96 = T655 & 32'hff00ff;
  assign T655 = {8'h0, T97};
  assign T97 = T89 >> 4'h8;
  assign T98 = T656 & 32'hf0f0f0f;
  assign T656 = {4'h0, T99};
  assign T99 = T85 >> 3'h4;
  assign T100 = T657 & 32'h33333333;
  assign T657 = {2'h0, T101};
  assign T101 = T81 >> 2'h2;
  assign T102 = T658 & 32'h55555555;
  assign T658 = {1'h0, T103};
  assign T103 = T77 >> 1'h1;
  assign T104 = 56'h0 - T659;
  assign T659 = {55'h0, T105};
  assign T105 = sExpX3[4'hd];
  assign sigX3 = T106[6'h38:1'h0];
  assign T106 = {T272, T107};
  assign T107 = doIncrSig ? T268 : T108;
  assign T108 = T109 != 32'h0;
  assign T109 = T178 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T110, 1'h1};
  assign T110 = {T153, T111};
  assign T111 = {T134, T112};
  assign T112 = {T124, T113};
  assign T113 = {T120, T114};
  assign T114 = T115[2'h2];
  assign T115 = T116[3'h6:3'h4];
  assign T116 = T117[4'he:4'h8];
  assign T117 = T118[5'h1e:5'h10];
  assign T118 = T119[5'h1f:1'h1];
  assign T119 = $signed(33'h100000000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = estNormDist[3'h4:1'h0];
  assign T120 = {T123, T121};
  assign T121 = T122[1'h1];
  assign T122 = T115[1'h1:1'h0];
  assign T123 = T122[1'h0];
  assign T124 = {T130, T125};
  assign T125 = {T129, T126};
  assign T126 = T127[1'h1];
  assign T127 = T128[2'h3:2'h2];
  assign T128 = T116[2'h3:1'h0];
  assign T129 = T127[1'h0];
  assign T130 = {T133, T131};
  assign T131 = T132[1'h1];
  assign T132 = T128[1'h1:1'h0];
  assign T133 = T132[1'h0];
  assign T134 = T151 | T135;
  assign T135 = T136 & 8'haa;
  assign T136 = T137 << 1'h1;
  assign T137 = T138[3'h6:1'h0];
  assign T138 = T149 | T139;
  assign T139 = T140 & 8'hcc;
  assign T140 = T141 << 2'h2;
  assign T141 = T142[3'h5:1'h0];
  assign T142 = T147 | T143;
  assign T143 = T144 & 8'hf0;
  assign T144 = T145 << 3'h4;
  assign T145 = T146[2'h3:1'h0];
  assign T146 = T117[3'h7:1'h0];
  assign T147 = T660 & 8'hf;
  assign T660 = {4'h0, T148};
  assign T148 = T146 >> 3'h4;
  assign T149 = T661 & 8'h33;
  assign T661 = {2'h0, T150};
  assign T150 = T142 >> 2'h2;
  assign T151 = T662 & 8'h55;
  assign T662 = {1'h0, T152};
  assign T152 = T138 >> 1'h1;
  assign T153 = T176 | T154;
  assign T154 = T155 & 16'haaaa;
  assign T155 = T156 << 1'h1;
  assign T156 = T157[4'he:1'h0];
  assign T157 = T174 | T158;
  assign T158 = T159 & 16'hcccc;
  assign T159 = T160 << 2'h2;
  assign T160 = T161[4'hd:1'h0];
  assign T161 = T172 | T162;
  assign T162 = T163 & 16'hf0f0;
  assign T163 = T164 << 3'h4;
  assign T164 = T165[4'hb:1'h0];
  assign T165 = T170 | T166;
  assign T166 = T167 & 16'hff00;
  assign T167 = T168 << 4'h8;
  assign T168 = T169[3'h7:1'h0];
  assign T169 = T118[4'hf:1'h0];
  assign T170 = T663 & 16'hff;
  assign T663 = {8'h0, T171};
  assign T171 = T169 >> 4'h8;
  assign T172 = T664 & 16'hf0f;
  assign T664 = {4'h0, T173};
  assign T173 = T165 >> 3'h4;
  assign T174 = T665 & 16'h3333;
  assign T665 = {2'h0, T175};
  assign T175 = T161 >> 2'h2;
  assign T176 = T666 & 16'h5555;
  assign T666 = {1'h0, T177};
  assign T177 = T157 >> 1'h1;
  assign T178 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T247 : T667;
  assign T667 = {1'h0, T179};
  assign T179 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T216 ? T204 : T180;
  assign T180 = T203 ? T184 : T181;
  assign T181 = {T183, T182};
  assign T182 = 54'h0 - T668;
  assign T668 = {53'h0, doSubMags};
  assign T183 = sigSum[6'h21:1'h1];
  assign T184 = T202 ? T670 : T185;
  assign T185 = {T187, T186};
  assign T186 = 86'h0 - T669;
  assign T669 = {85'h0, doSubMags};
  assign T187 = sigSum[1'h1];
  assign T670 = {21'h0, T188};
  assign T188 = {T201, T189};
  assign T189 = doSubMags ? T195 : T190;
  assign T190 = firstReduceSigSum[1'h0];
  assign firstReduceSigSum = {T193, T191};
  assign T191 = T192 != 44'h0;
  assign T192 = sigSum[6'h2b:1'h0];
  assign T193 = T194 != 32'h0;
  assign T194 = sigSum[7'h4b:6'h2c];
  assign T195 = T196 ^ 1'h1;
  assign T196 = firstReduceComplSigSum[1'h0];
  assign firstReduceComplSigSum = {T199, T197};
  assign T197 = T198 != 44'h0;
  assign T198 = complSigSum[6'h2b:1'h0];
  assign complSigSum = ~ sigSum;
  assign T199 = T200 != 32'h0;
  assign T200 = complSigSum[7'h4b:6'h2c];
  assign T201 = sigSum[7'h6c:6'h2c];
  assign T202 = estNormNeg_dist[3'h4];
  assign T203 = estNormNeg_dist[3'h5];
  assign T204 = T215 ? T212 : T205;
  assign T205 = {T211, T206};
  assign T206 = doSubMags ? T209 : T207;
  assign T207 = T208 != 11'h0;
  assign T208 = sigSum[4'hb:1'h1];
  assign T209 = T210 == 11'h0;
  assign T210 = complSigSum[4'hb:1'h1];
  assign T211 = sigSum[7'h61:4'hc];
  assign T212 = {T214, T213};
  assign T213 = 22'h0 - T671;
  assign T671 = {21'h0, doSubMags};
  assign T214 = sigSum[7'h41:1'h1];
  assign T215 = estNormNeg_dist[3'h5];
  assign T216 = estNormNeg_dist[3'h6];
  assign CDom_firstNormAbsSigSum = T223 | T217;
  assign T217 = T221 ? T218 : 87'h0;
  assign T218 = {T220, T219};
  assign T219 = firstReduceComplSigSum[1'h0];
  assign T220 = complSigSum[8'h81:6'h2c];
  assign T221 = doSubMags & T222;
  assign T222 = CDom_estNormDist[3'h5];
  assign T223 = T231 | T224;
  assign T224 = T228 ? T225 : 87'h0;
  assign T225 = {T227, T226};
  assign T226 = firstReduceComplSigSum != 2'h0;
  assign T227 = complSigSum[8'ha1:7'h4c];
  assign T228 = doSubMags & T229;
  assign T229 = T230 ^ 1'h1;
  assign T230 = CDom_estNormDist[3'h5];
  assign T231 = T239 | T232;
  assign T232 = T236 ? T233 : 87'h0;
  assign T233 = {T235, T234};
  assign T234 = firstReduceSigSum[1'h0];
  assign T235 = sigSum[8'h81:6'h2c];
  assign T236 = T238 & T237;
  assign T237 = CDom_estNormDist[3'h5];
  assign T238 = doSubMags ^ 1'h1;
  assign T239 = T243 ? T240 : 87'h0;
  assign T240 = {T242, T241};
  assign T241 = firstReduceSigSum != 2'h0;
  assign T242 = sigSum[8'ha1:7'h4c];
  assign T243 = T246 & T244;
  assign T244 = T245 ^ 1'h1;
  assign T245 = CDom_estNormDist[3'h5];
  assign T246 = doSubMags ^ 1'h1;
  assign T247 = io_fromPreMul_isCDominant ? T673 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T267 ? T259 : T248;
  assign T248 = T258 ? T251 : T249;
  assign T249 = T250 << 6'h36;
  assign T250 = complSigSum[6'h22:1'h1];
  assign T251 = T257 ? T672 : T252;
  assign T252 = T253 << 7'h56;
  assign T253 = complSigSum[2'h2:1'h1];
  assign T672 = {23'h0, T254};
  assign T254 = {T256, T255};
  assign T255 = firstReduceComplSigSum[1'h0];
  assign T256 = complSigSum[7'h6b:6'h2c];
  assign T257 = estNormNeg_dist[3'h4];
  assign T258 = estNormNeg_dist[3'h5];
  assign T259 = T266 ? T264 : T260;
  assign T260 = {T263, T261};
  assign T261 = T262 != 11'h0;
  assign T262 = complSigSum[4'hb:1'h1];
  assign T263 = complSigSum[7'h62:4'hc];
  assign T264 = T265 << 5'h16;
  assign T265 = complSigSum[7'h42:1'h1];
  assign T266 = estNormNeg_dist[3'h5];
  assign T267 = estNormNeg_dist[3'h6];
  assign T673 = {1'h0, CDom_firstNormAbsSigSum};
  assign T268 = T269 == 32'h0;
  assign T269 = T270 & absSigSumExtraMask;
  assign T270 = ~ T271;
  assign T271 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign T272 = T273 >> normTo2ShiftDist;
  assign T273 = cFirstNormAbsSigSum[7'h57:1'h1];
  assign roundPosBit = T274 != 57'h0;
  assign T274 = sigX3 & T674;
  assign T674 = {1'h0, roundPosMask};
  assign roundPosMask = T675 & roundMask;
  assign T675 = {1'h0, T275};
  assign T275 = ~ T276;
  assign T276 = roundMask >> 1'h1;
  assign T277 = allRound ^ 1'h1;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T278 == 57'h0;
  assign T278 = T280 & T676;
  assign T676 = {2'h0, T279};
  assign T279 = roundMask >> 1'h1;
  assign T280 = ~ sigX3;
  assign doIncrSig = T281 & doSubMags;
  assign T281 = T283 & T282;
  assign T282 = notCDom_signSigSum ^ 1'h1;
  assign T283 = io_fromPreMul_isCDominant ^ 1'h1;
  assign commonCase = T285 & T284;
  assign T284 = notSpecial_addZeros ^ 1'h1;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign isZeroC = io_fromPreMul_highExpC == 3'h0;
  assign T285 = addSpecial ^ 1'h1;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T286 == 2'h3;
  assign T286 = io_fromPreMul_highExpC[2'h2:1'h1];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T287 == 2'h3;
  assign T287 = io_fromPreMul_highExpB[2'h2:1'h1];
  assign isSpecialA = T288 == 2'h3;
  assign T288 = io_fromPreMul_highExpA[2'h2:1'h1];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T289;
  assign T289 = T293 | T290;
  assign T290 = sExpX3_13 <= T677;
  assign T677 = {2'h0, T291};
  assign T291 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign sigX3Shift1 = T292 == 2'h0;
  assign T292 = sigX3[6'h38:6'h37];
  assign T293 = sExpX3[4'hd];
  assign overflow = commonCase & overflowY;
  assign overflowY = T294 == 3'h3;
  assign T294 = sExpY[4'hc:4'ha];
  assign sExpY = T339 | T295;
  assign T295 = T297 ? T296 : 14'h0;
  assign T296 = sExpX3 - 14'h1;
  assign T297 = T298 == 2'h0;
  assign T298 = sigY3[6'h36:6'h35];
  assign sigY3 = T312 | T299;
  assign T299 = roundEven ? T300 : 55'h0;
  assign T300 = roundUp_sigY3 & T301;
  assign T301 = ~ T302;
  assign T302 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T303;
  assign T303 = T304 + 55'h1;
  assign T304 = T305 >> 2'h2;
  assign T305 = sigX3 | T678;
  assign T678 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T309 : T306;
  assign T306 = T308 & T307;
  assign T307 = anyRoundExtra ^ 1'h1;
  assign T308 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign T309 = T310 & allRoundExtra;
  assign T310 = roundingMode_nearest_even & T311;
  assign T311 = roundPosBit ^ 1'h1;
  assign T312 = T332 | T313;
  assign T313 = roundUp ? roundUp_sigY3 : 55'h0;
  assign roundUp = T319 | T314;
  assign T314 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign signY = isZeroY ? roundingMode_min : T315;
  assign T315 = io_fromPreMul_signProd ^ doNegSignSum;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T316 : notCDom_signSigSum;
  assign T316 = doSubMags & T317;
  assign T317 = isZeroC ^ 1'h1;
  assign isZeroY = T318 == 3'h0;
  assign T318 = sigX3[6'h38:6'h36];
  assign T319 = T322 | T320;
  assign T320 = T321 & roundPosBit;
  assign T321 = doIncrSig & roundingMode_nearest_even;
  assign T322 = T324 | T323;
  assign T323 = doIncrSig & allRound;
  assign T324 = T328 | T325;
  assign T325 = T326 & anyRound;
  assign T326 = T327 & roundDirectUp;
  assign T327 = doIncrSig ^ 1'h1;
  assign T328 = T329 & anyRoundExtra;
  assign T329 = T330 & roundPosBit;
  assign T330 = T331 & roundingMode_nearest_even;
  assign T331 = doIncrSig ^ 1'h1;
  assign T332 = T336 ? T333 : 55'h0;
  assign T333 = T334 >> 2'h2;
  assign T334 = sigX3 & T679;
  assign T679 = {1'h0, T335};
  assign T335 = ~ roundMask;
  assign T336 = T338 & T337;
  assign T337 = roundEven ^ 1'h1;
  assign T338 = roundUp ^ 1'h1;
  assign T339 = T342 | T340;
  assign T340 = T341 ? sExpX3 : 14'h0;
  assign T341 = sigY3[6'h35];
  assign T342 = T344 ? T343 : 14'h0;
  assign T343 = sExpX3 + 14'h1;
  assign T344 = sigY3[6'h36];
  assign T345 = {invalid, 1'h0};
  assign invalid = T364 | notSigNaN_invalid;
  assign notSigNaN_invalid = T361 | T346;
  assign T346 = T347 & doSubMags;
  assign T347 = T350 & isInfC;
  assign isInfC = isSpecialC & T348;
  assign T348 = T349 ^ 1'h1;
  assign T349 = io_fromPreMul_highExpC[1'h0];
  assign T350 = T356 & T351;
  assign T351 = isInfA | isInfB;
  assign isInfB = isSpecialB & T352;
  assign T352 = T353 ^ 1'h1;
  assign T353 = io_fromPreMul_highExpB[1'h0];
  assign isInfA = isSpecialA & T354;
  assign T354 = T355 ^ 1'h1;
  assign T355 = io_fromPreMul_highExpA[1'h0];
  assign T356 = T359 & T357;
  assign T357 = isNaNB ^ 1'h1;
  assign isNaNB = isSpecialB & T358;
  assign T358 = io_fromPreMul_highExpB[1'h0];
  assign T359 = isNaNA ^ 1'h1;
  assign isNaNA = isSpecialA & T360;
  assign T360 = io_fromPreMul_highExpA[1'h0];
  assign T361 = T363 | T362;
  assign T362 = isZeroA & isInfB;
  assign isZeroA = io_fromPreMul_highExpA == 3'h0;
  assign T363 = isInfA & isZeroB;
  assign isZeroB = io_fromPreMul_highExpB == 3'h0;
  assign T364 = T367 | isSigNaNC;
  assign isSigNaNC = isNaNC & T365;
  assign T365 = io_fromPreMul_isNaN_isQuietNaNC ^ 1'h1;
  assign isNaNC = isSpecialC & T366;
  assign T366 = io_fromPreMul_highExpC[1'h0];
  assign T367 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T368;
  assign T368 = io_fromPreMul_isNaN_isQuietNaNB ^ 1'h1;
  assign isSigNaNA = isNaNA & T369;
  assign T369 = io_fromPreMul_isNaN_isQuietNaNA ^ 1'h1;
  assign io_out = T370;
  assign T370 = {signOut, T371};
  assign T371 = {expOut, fractOut};
  assign fractOut = T377 | T372;
  assign T372 = 52'h0 - T680;
  assign T680 = {51'h0, pegMaxFiniteMagOut};
  assign pegMaxFiniteMagOut = overflow & T373;
  assign T373 = overflowY_roundMagUp ^ 1'h1;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign roundMagUp = T376 | T374;
  assign T374 = roundingMode_max & T375;
  assign T375 = signY ^ 1'h1;
  assign T376 = roundingMode_min & signY;
  assign T377 = T383 ? T380 : fractY;
  assign fractY = sigX3Shift1 ? T379 : T378;
  assign T378 = sigY3[6'h34:1'h1];
  assign T379 = sigY3[6'h33:1'h0];
  assign T380 = isNaNOut ? 52'h8000000000000 : 52'h0;
  assign isNaNOut = T381 | notSigNaN_invalid;
  assign T381 = T382 | isNaNC;
  assign T382 = isNaNA | isNaNB;
  assign T383 = T384 | isNaNOut;
  assign T384 = totalUnderflowY & roundMagUp;
  assign totalUnderflowY = T389 & T385;
  assign T385 = T388 | T386;
  assign T386 = T387 < 12'h3ce;
  assign T387 = sExpY[4'hb:1'h0];
  assign T388 = sExpY[4'hc];
  assign T389 = isZeroY ^ 1'h1;
  assign expOut = T391 | T390;
  assign T390 = isNaNOut ? 12'he00 : 12'h0;
  assign T391 = T396 | T392;
  assign T392 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = T394 | T393;
  assign T393 = overflow & overflowY_roundMagUp;
  assign T394 = T395 | isInfC;
  assign T395 = isInfA | isInfB;
  assign T396 = T398 | T397;
  assign T397 = pegMaxFiniteMagOut ? 12'hbff : 12'h0;
  assign T398 = T401 | T399;
  assign T399 = pegMinFiniteMagOut ? 12'h3ce : 12'h0;
  assign pegMinFiniteMagOut = T400 & roundMagUp;
  assign T400 = commonCase & totalUnderflowY;
  assign T401 = T404 & T402;
  assign T402 = ~ T403;
  assign T403 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T404 = T407 & T405;
  assign T405 = ~ T406;
  assign T406 = pegMaxFiniteMagOut ? 12'h400 : 12'h0;
  assign T407 = T410 & T408;
  assign T408 = ~ T409;
  assign T409 = pegMinFiniteMagOut ? 12'hc31 : 12'h0;
  assign T410 = expY & T411;
  assign T411 = ~ T412;
  assign T412 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign notSpecial_isZeroOut = T413 | totalUnderflowY;
  assign T413 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'hb:1'h0];
  assign signOut = T415 | T414;
  assign T414 = commonCase & signY;
  assign T415 = T430 & uncommonCaseSignOut;
  assign uncommonCaseSignOut = T420 | T416;
  assign T416 = T417 & roundingMode_min;
  assign T417 = T418 & doSubMags;
  assign T418 = T419 & notSpecial_addZeros;
  assign T419 = mulSpecial ^ 1'h1;
  assign T420 = T424 | T421;
  assign T421 = T422 & io_fromPreMul_opSignC;
  assign T422 = T423 & isSpecialC;
  assign T423 = mulSpecial ^ 1'h1;
  assign T424 = T428 | T425;
  assign T425 = T426 & io_fromPreMul_signProd;
  assign T426 = mulSpecial & T427;
  assign T427 = isSpecialC ^ 1'h1;
  assign T428 = T429 & io_fromPreMul_opSignC;
  assign T429 = doSubMags ^ 1'h1;
  assign T430 = isNaNOut ^ 1'h1;
endmodule

module MulAddRecFN_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[106:0] T0;
  wire[106:0] T1;
  wire[106:0] T3;
  wire[105:0] T2;
  wire[52:0] mulAddRecFN_preMul_io_mulAddA;
  wire[52:0] mulAddRecFN_preMul_io_mulAddB;
  wire[105:0] mulAddRecFN_preMul_io_mulAddC;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire mulAddRecFN_preMul_io_toPostMul_signProd;
  wire mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire[2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire[7:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire[54:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire[13:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire[1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire[64:0] mulAddRecFN_postMul_io_out;
  wire[4:0] mulAddRecFN_postMul_io_exceptionFlags;


  assign T0 = T3 + T1;
  assign T1 = {1'h0, mulAddRecFN_preMul_io_mulAddC};
  assign T3 = {1'h0, T2};
  assign T2 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign io_out = mulAddRecFN_postMul_io_out;
  MulAddRecFN_preMul_1 mulAddRecFN_preMul(
       .io_op( io_op ),
       .io_a( io_a ),
       .io_b( io_b ),
       .io_c( io_c ),
       .io_roundingMode( io_roundingMode ),
       .io_mulAddA( mulAddRecFN_preMul_io_mulAddA ),
       .io_mulAddB( mulAddRecFN_preMul_io_mulAddB ),
       .io_mulAddC( mulAddRecFN_preMul_io_mulAddC ),
       .io_toPostMul_highExpA( mulAddRecFN_preMul_io_toPostMul_highExpA ),
       .io_toPostMul_isNaN_isQuietNaNA( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA ),
       .io_toPostMul_highExpB( mulAddRecFN_preMul_io_toPostMul_highExpB ),
       .io_toPostMul_isNaN_isQuietNaNB( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB ),
       .io_toPostMul_signProd( mulAddRecFN_preMul_io_toPostMul_signProd ),
       .io_toPostMul_isZeroProd( mulAddRecFN_preMul_io_toPostMul_isZeroProd ),
       .io_toPostMul_opSignC( mulAddRecFN_preMul_io_toPostMul_opSignC ),
       .io_toPostMul_highExpC( mulAddRecFN_preMul_io_toPostMul_highExpC ),
       .io_toPostMul_isNaN_isQuietNaNC( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC ),
       .io_toPostMul_isCDominant( mulAddRecFN_preMul_io_toPostMul_isCDominant ),
       .io_toPostMul_CAlignDist_0( mulAddRecFN_preMul_io_toPostMul_CAlignDist_0 ),
       .io_toPostMul_CAlignDist( mulAddRecFN_preMul_io_toPostMul_CAlignDist ),
       .io_toPostMul_bit0AlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC ),
       .io_toPostMul_highAlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC ),
       .io_toPostMul_sExpSum( mulAddRecFN_preMul_io_toPostMul_sExpSum ),
       .io_toPostMul_roundingMode( mulAddRecFN_preMul_io_toPostMul_roundingMode )
  );
  MulAddRecFN_postMul_1 mulAddRecFN_postMul(
       .io_fromPreMul_highExpA( mulAddRecFN_preMul_io_toPostMul_highExpA ),
       .io_fromPreMul_isNaN_isQuietNaNA( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA ),
       .io_fromPreMul_highExpB( mulAddRecFN_preMul_io_toPostMul_highExpB ),
       .io_fromPreMul_isNaN_isQuietNaNB( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB ),
       .io_fromPreMul_signProd( mulAddRecFN_preMul_io_toPostMul_signProd ),
       .io_fromPreMul_isZeroProd( mulAddRecFN_preMul_io_toPostMul_isZeroProd ),
       .io_fromPreMul_opSignC( mulAddRecFN_preMul_io_toPostMul_opSignC ),
       .io_fromPreMul_highExpC( mulAddRecFN_preMul_io_toPostMul_highExpC ),
       .io_fromPreMul_isNaN_isQuietNaNC( mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC ),
       .io_fromPreMul_isCDominant( mulAddRecFN_preMul_io_toPostMul_isCDominant ),
       .io_fromPreMul_CAlignDist_0( mulAddRecFN_preMul_io_toPostMul_CAlignDist_0 ),
       .io_fromPreMul_CAlignDist( mulAddRecFN_preMul_io_toPostMul_CAlignDist ),
       .io_fromPreMul_bit0AlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC ),
       .io_fromPreMul_highAlignedNegSigC( mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC ),
       .io_fromPreMul_sExpSum( mulAddRecFN_preMul_io_toPostMul_sExpSum ),
       .io_fromPreMul_roundingMode( mulAddRecFN_preMul_io_toPostMul_roundingMode ),
       .io_mulAddResult( T0 ),
       .io_out( mulAddRecFN_postMul_io_out ),
       .io_exceptionFlags( mulAddRecFN_postMul_io_exceptionFlags )
  );
endmodule

module FPUFMAPipe_1(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap12,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_div,
    input  io_in_bits_sqrt,
    input  io_in_bits_round,
    input  io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T31;
  reg [2:0] in_rm;
  wire[2:0] T0;
  reg [64:0] in_in3;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[64:0] zero;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] in_in2;
  wire[64:0] T9;
  wire[64:0] T10;
  wire T11;
  reg [64:0] in_in1;
  wire[64:0] T12;
  wire[1:0] T32;
  reg [4:0] in_cmd;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T33;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [4:0] R20;
  wire[4:0] T21;
  reg [4:0] R22;
  wire[4:0] T23;
  wire[4:0] res_exc;
  reg  valid;
  reg  R24;
  wire T34;
  reg [64:0] R25;
  wire[64:0] T26;
  reg [64:0] R27;
  wire[64:0] T28;
  wire[64:0] res_data;
  wire[64:0] T35;
  wire[96:0] T29;
  reg  R30;
  wire T36;
  wire[64:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R20 = {1{$random}};
    R22 = {1{$random}};
    valid = {1{$random}};
    R24 = {1{$random}};
    R25 = {3{$random}};
    R27 = {3{$random}};
    R30 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T31 = in_rm[1'h1:1'h0];
  assign T0 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T1 = T6 ? zero : T2;
  assign T2 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign zero = T3 << 7'h40;
  assign T3 = T5 ^ T4;
  assign T4 = io_in_bits_in2[7'h40];
  assign T5 = io_in_bits_in1[7'h40];
  assign T6 = io_in_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T9 = T11 ? 65'h8000000000000000 : T10;
  assign T10 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T11 = io_in_valid & io_in_bits_swap23;
  assign T12 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T32 = in_cmd[1'h1:1'h0];
  assign T13 = io_in_valid ? T33 : T14;
  assign T14 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T33 = {3'h0, T15};
  assign T15 = {T17, T16};
  assign T16 = io_in_bits_cmd[1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = io_in_bits_cmd[1'h1];
  assign io_out_bits_exc = R20;
  assign T21 = R24 ? R22 : R20;
  assign T23 = valid ? res_exc : R22;
  assign res_exc = fma_io_exceptionFlags;
  assign T34 = reset ? 1'h0 : valid;
  assign io_out_bits_data = R25;
  assign T26 = R24 ? R27 : R25;
  assign T28 = valid ? res_data : R27;
  assign res_data = T35;
  assign T35 = T29[7'h40:1'h0];
  assign T29 = {32'hffffffff, fma_io_out};
  assign io_out_valid = R30;
  assign T36 = reset ? 1'h0 : R24;
  MulAddRecFN_1 fma(
       .io_op( T32 ),
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_c( in_in3 ),
       .io_roundingMode( T31 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T6) begin
      in_in3 <= zero;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T11) begin
      in_in2 <= 65'h8000000000000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T33;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(R24) begin
      R20 <= R22;
    end
    if(valid) begin
      R22 <= res_exc;
    end
    valid <= io_in_valid;
    if(reset) begin
      R24 <= 1'h0;
    end else begin
      R24 <= valid;
    end
    if(R24) begin
      R25 <= R27;
    end
    if(valid) begin
      R27 <= res_data;
    end
    if(reset) begin
      R30 <= 1'h0;
    end else begin
      R30 <= R24;
    end
  end
endmodule

module RecFNToRecFN(
    input [32:0] io_in,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire invalidExc;
  wire T1;
  wire T2;
  wire[55:0] outRawFloat_sig;
  wire[55:0] T3;
  wire[26:0] T4;
  wire[26:0] T5;
  wire[24:0] T6;
  wire[22:0] T7;
  wire outRawFloat_isNaN;
  wire T8;
  wire T9;
  wire T10;
  wire[8:0] T11;
  wire T12;
  wire[1:0] T13;
  wire[64:0] T14;
  wire[63:0] T15;
  wire[51:0] T16;
  wire[51:0] T17;
  wire[11:0] T18;
  wire[11:0] T19;
  wire[11:0] T20;
  wire[11:0] T21;
  wire outRawFloat_isInf;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[11:0] T26;
  wire[11:0] T27;
  wire[11:0] T28;
  wire T29;
  wire outRawFloat_isZero;
  wire T30;
  wire T31;
  wire[2:0] T32;
  wire[11:0] T33;
  wire[11:0] T34;
  wire[11:0] T35;
  wire[11:0] T36;
  wire[12:0] outRawFloat_sExp;
  wire[12:0] T45;
  wire[11:0] T37;
  wire[11:0] T46;
  wire[9:0] T38;
  wire[9:0] T39;
  wire[9:0] T40;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T41;
  wire T42;
  wire outRawFloat_sign;
  wire T43;
  wire T44;


  assign io_exceptionFlags = T0;
  assign T0 = {invalidExc, 4'h0};
  assign invalidExc = outRawFloat_isNaN & T1;
  assign T1 = T2 ^ 1'h1;
  assign T2 = outRawFloat_sig[6'h35];
  assign outRawFloat_sig = T3;
  assign T3 = T4 << 5'h1d;
  assign T4 = T5;
  assign T5 = {2'h1, T6};
  assign T6 = {T7, 2'h0};
  assign T7 = io_in[5'h16:1'h0];
  assign outRawFloat_isNaN = T8;
  assign T8 = T9;
  assign T9 = T12 & T10;
  assign T10 = T11[3'h6];
  assign T11 = io_in[5'h1f:5'h17];
  assign T12 = T13 == 2'h3;
  assign T13 = T11[4'h8:3'h7];
  assign io_out = T14;
  assign T14 = {T41, T15};
  assign T15 = {T18, T16};
  assign T16 = outRawFloat_isNaN ? 52'h8000000000000 : T17;
  assign T17 = outRawFloat_sig[6'h35:2'h2];
  assign T18 = T20 | T19;
  assign T19 = outRawFloat_isNaN ? 12'he00 : 12'h0;
  assign T20 = T26 | T21;
  assign T21 = outRawFloat_isInf ? 12'hc00 : 12'h0;
  assign outRawFloat_isInf = T22;
  assign T22 = T23;
  assign T23 = T12 & T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = T11[3'h6];
  assign T26 = T33 & T27;
  assign T27 = ~ T28;
  assign T28 = T29 ? 12'h200 : 12'h0;
  assign T29 = outRawFloat_isZero | outRawFloat_isInf;
  assign outRawFloat_isZero = T30;
  assign T30 = T31;
  assign T31 = T32 == 3'h0;
  assign T32 = T11[4'h8:3'h6];
  assign T33 = T36 & T34;
  assign T34 = ~ T35;
  assign T35 = outRawFloat_isZero ? 12'hc00 : 12'h0;
  assign T36 = outRawFloat_sExp[4'hb:1'h0];
  assign outRawFloat_sExp = T45;
  assign T45 = {T49, T37};
  assign T37 = T46 + 12'h700;
  assign T46 = {T47, T38};
  assign T38 = T39;
  assign T39 = T40;
  assign T40 = {1'h0, T11};
  assign T47 = T48 ? 2'h3 : 2'h0;
  assign T48 = T38[4'h9];
  assign T49 = T37[4'hb];
  assign T41 = outRawFloat_sign & T42;
  assign T42 = outRawFloat_isNaN ^ 1'h1;
  assign outRawFloat_sign = T43;
  assign T43 = T44;
  assign T44 = io_in[6'h20];
endmodule

module CompareRecFN(
    input [64:0] io_a,
    input [64:0] io_b,
    input  io_signaling,
    output io_lt,
    output io_eq,
    output io_gt,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire invalid;
  wire T1;
  wire T2;
  wire ordered;
  wire T3;
  wire rawB_isNaN;
  wire T4;
  wire T5;
  wire[11:0] T6;
  wire T7;
  wire[1:0] T8;
  wire T9;
  wire rawA_isNaN;
  wire T10;
  wire T11;
  wire[11:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[55:0] rawB_sig;
  wire[55:0] T19;
  wire[53:0] T20;
  wire[51:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[55:0] rawA_sig;
  wire[55:0] T25;
  wire[53:0] T26;
  wire[51:0] T27;
  wire T28;
  wire T29;
  wire ordered_eq;
  wire T30;
  wire T31;
  wire common_eqMags;
  wire T32;
  wire eqExps;
  wire[12:0] rawB_sExp;
  wire[12:0] T33;
  wire[12:0] T34;
  wire[12:0] rawA_sExp;
  wire[12:0] T35;
  wire[12:0] T36;
  wire bothInfs;
  wire rawB_isInf;
  wire T37;
  wire T38;
  wire T39;
  wire rawA_isInf;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire rawB_sign;
  wire T44;
  wire rawA_sign;
  wire T45;
  wire bothZeros;
  wire rawB_isZero;
  wire T46;
  wire[2:0] T47;
  wire rawA_isZero;
  wire T48;
  wire[2:0] T49;
  wire T50;
  wire T51;
  wire ordered_lt;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire common_ltMags;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;


  assign io_exceptionFlags = T0;
  assign T0 = {invalid, 4'h0};
  assign invalid = T15 | T1;
  assign T1 = io_signaling & T2;
  assign T2 = ordered ^ 1'h1;
  assign ordered = T9 & T3;
  assign T3 = rawB_isNaN ^ 1'h1;
  assign rawB_isNaN = T4;
  assign T4 = T7 & T5;
  assign T5 = T6[4'h9];
  assign T6 = io_b[6'h3f:6'h34];
  assign T7 = T8 == 2'h3;
  assign T8 = T6[4'hb:4'ha];
  assign T9 = rawA_isNaN ^ 1'h1;
  assign rawA_isNaN = T10;
  assign T10 = T13 & T11;
  assign T11 = T12[4'h9];
  assign T12 = io_a[6'h3f:6'h34];
  assign T13 = T14 == 2'h3;
  assign T14 = T12[4'hb:4'ha];
  assign T15 = T22 | T16;
  assign T16 = rawB_isNaN & T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = rawB_sig[6'h35];
  assign rawB_sig = T19;
  assign T19 = {2'h1, T20};
  assign T20 = {T21, 2'h0};
  assign T21 = io_b[6'h33:1'h0];
  assign T22 = rawA_isNaN & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = rawA_sig[6'h35];
  assign rawA_sig = T25;
  assign T25 = {2'h1, T26};
  assign T26 = {T27, 2'h0};
  assign T27 = io_a[6'h33:1'h0];
  assign io_gt = T28;
  assign T28 = T50 & T29;
  assign T29 = ordered_eq ^ 1'h1;
  assign ordered_eq = bothZeros | T30;
  assign T30 = T43 & T31;
  assign T31 = bothInfs | common_eqMags;
  assign common_eqMags = eqExps & T32;
  assign T32 = rawA_sig == rawB_sig;
  assign eqExps = rawA_sExp == rawB_sExp;
  assign rawB_sExp = T33;
  assign T33 = T34;
  assign T34 = {1'h0, T6};
  assign rawA_sExp = T35;
  assign T35 = T36;
  assign T36 = {1'h0, T12};
  assign bothInfs = rawA_isInf & rawB_isInf;
  assign rawB_isInf = T37;
  assign T37 = T7 & T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T6[4'h9];
  assign rawA_isInf = T40;
  assign T40 = T13 & T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T12[4'h9];
  assign T43 = rawA_sign == rawB_sign;
  assign rawB_sign = T44;
  assign T44 = io_b[7'h40];
  assign rawA_sign = T45;
  assign T45 = io_a[7'h40];
  assign bothZeros = rawA_isZero & rawB_isZero;
  assign rawB_isZero = T46;
  assign T46 = T47 == 3'h0;
  assign T47 = T6[4'hb:4'h9];
  assign rawA_isZero = T48;
  assign T48 = T49 == 3'h0;
  assign T49 = T12[4'hb:4'h9];
  assign T50 = ordered & T51;
  assign T51 = ordered_lt ^ 1'h1;
  assign ordered_lt = T67 & T52;
  assign T52 = T65 | T53;
  assign T53 = T64 & T54;
  assign T54 = T60 | T55;
  assign T55 = T59 & common_ltMags;
  assign common_ltMags = T58 | T56;
  assign T56 = eqExps & T57;
  assign T57 = rawA_sig < rawB_sig;
  assign T58 = $signed(rawA_sExp) < $signed(rawB_sExp);
  assign T59 = rawB_sign ^ 1'h1;
  assign T60 = T62 & T61;
  assign T61 = common_eqMags ^ 1'h1;
  assign T62 = rawA_sign & T63;
  assign T63 = common_ltMags ^ 1'h1;
  assign T64 = bothInfs ^ 1'h1;
  assign T65 = rawA_sign & T66;
  assign T66 = rawB_sign ^ 1'h1;
  assign T67 = bothZeros ^ 1'h1;
  assign io_eq = T68;
  assign T68 = ordered & ordered_eq;
  assign io_lt = T69;
  assign T69 = ordered & ordered_lt;
endmodule

module RecFNToIN_0(
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    input  io_signedOut,
    output[63:0] io_out,
    output[2:0] io_intExceptionFlags
);

  wire[2:0] T0;
  wire[1:0] T1;
  wire inexact;
  wire T2;
  wire T3;
  wire T4;
  wire roundInexact;
  wire T5;
  wire isZero;
  wire[2:0] T6;
  wire[11:0] exp;
  wire T7;
  wire[1:0] T8;
  wire[2:0] roundBits;
  wire T9;
  wire[50:0] T10;
  wire[115:0] shiftedSig;
  wire[5:0] T11;
  wire[5:0] T12;
  wire[52:0] T13;
  wire[51:0] fract;
  wire[1:0] T14;
  wire notSpecial_magGeOne;
  wire overflow;
  wire overflow_unsigned;
  wire T15;
  wire roundIncr;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire roundIncr_nearestEven;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire T28;
  wire[10:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire sign;
  wire T36;
  wire T37;
  wire roundCarryBut2;
  wire T38;
  wire[61:0] T39;
  wire[63:0] unroundedInt;
  wire T40;
  wire T41;
  wire T42;
  wire[10:0] posExp;
  wire T43;
  wire T44;
  wire overflow_signed;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[62:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire invalid;
  wire[1:0] T59;
  wire[63:0] T60;
  wire[63:0] roundedInt;
  wire[63:0] complUnroundedInt;
  wire[63:0] T61;
  wire[63:0] T62;
  wire T63;
  wire[63:0] excValue;
  wire[63:0] T64;
  wire T65;
  wire T66;
  wire excSign;
  wire T67;
  wire isNaN;
  wire T68;
  wire T69;
  wire[63:0] T70;
  wire[63:0] T77;
  wire[62:0] T71;
  wire T72;
  wire T73;
  wire[63:0] T74;
  wire T75;
  wire T76;


  assign io_intExceptionFlags = T0;
  assign T0 = {invalid, T1};
  assign T1 = {overflow, inexact};
  assign inexact = T3 & T2;
  assign T2 = overflow ^ 1'h1;
  assign T3 = roundInexact & T4;
  assign T4 = invalid ^ 1'h1;
  assign roundInexact = notSpecial_magGeOne ? T7 : T5;
  assign T5 = isZero ^ 1'h1;
  assign isZero = T6 == 3'h0;
  assign T6 = exp[4'hb:4'h9];
  assign exp = io_in[6'h3f:6'h34];
  assign T7 = T8 != 2'h0;
  assign T8 = roundBits[1'h1:1'h0];
  assign roundBits = {T14, T9};
  assign T9 = T10 != 51'h0;
  assign T10 = shiftedSig[6'h32:1'h0];
  assign shiftedSig = T13 << T11;
  assign T11 = notSpecial_magGeOne ? T12 : 6'h0;
  assign T12 = exp[3'h5:1'h0];
  assign T13 = {notSpecial_magGeOne, fract};
  assign fract = io_in[6'h33:1'h0];
  assign T14 = shiftedSig[6'h34:6'h33];
  assign notSpecial_magGeOne = exp[4'hb];
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign overflow_unsigned = notSpecial_magGeOne ? T36 : T15;
  assign T15 = sign & roundIncr;
  assign roundIncr = T20 | T16;
  assign T16 = T19 & T17;
  assign T17 = T18 & roundInexact;
  assign T18 = sign ^ 1'h1;
  assign T19 = io_roundingMode == 2'h3;
  assign T20 = T24 | T21;
  assign T21 = T23 & T22;
  assign T22 = sign & roundInexact;
  assign T23 = io_roundingMode == 2'h2;
  assign T24 = T35 & roundIncr_nearestEven;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T30 : T25;
  assign T25 = T28 ? T26 : 1'h0;
  assign T26 = T27 != 2'h0;
  assign T27 = roundBits[1'h1:1'h0];
  assign T28 = T29 == 11'h7ff;
  assign T29 = exp[4'ha:1'h0];
  assign T30 = T33 | T31;
  assign T31 = T32 == 2'h3;
  assign T32 = roundBits[1'h1:1'h0];
  assign T33 = T34 == 2'h3;
  assign T34 = roundBits[2'h2:1'h1];
  assign T35 = io_roundingMode == 2'h0;
  assign sign = io_in[7'h40];
  assign T36 = T43 | T37;
  assign T37 = T40 & roundCarryBut2;
  assign roundCarryBut2 = T38 & roundIncr;
  assign T38 = T39 == 62'h3fffffffffffffff;
  assign T39 = unroundedInt[6'h3d:1'h0];
  assign unroundedInt = shiftedSig[7'h73:6'h34];
  assign T40 = T42 & T41;
  assign T41 = unroundedInt[6'h3e];
  assign T42 = posExp == 11'h3f;
  assign posExp = exp[4'ha:1'h0];
  assign T43 = sign | T44;
  assign T44 = 11'h40 <= posExp;
  assign overflow_signed = notSpecial_magGeOne ? T45 : 1'h0;
  assign T45 = T50 | T46;
  assign T46 = T47 & roundCarryBut2;
  assign T47 = T49 & T48;
  assign T48 = posExp == 11'h3e;
  assign T49 = sign ^ 1'h1;
  assign T50 = T58 | T51;
  assign T51 = T57 & T52;
  assign T52 = T53 | roundIncr;
  assign T53 = T56 | T54;
  assign T54 = T55 != 63'h0;
  assign T55 = unroundedInt[6'h3e:1'h0];
  assign T56 = sign ^ 1'h1;
  assign T57 = posExp == 11'h3f;
  assign T58 = 11'h40 <= posExp;
  assign invalid = T59 == 2'h3;
  assign T59 = exp[4'hb:4'ha];
  assign io_out = T60;
  assign T60 = T76 ? excValue : roundedInt;
  assign roundedInt = T63 ? T62 : complUnroundedInt;
  assign complUnroundedInt = sign ? T61 : unroundedInt;
  assign T61 = ~ unroundedInt;
  assign T62 = complUnroundedInt + 64'h1;
  assign T63 = roundIncr ^ sign;
  assign excValue = T70 | T64;
  assign T64 = T65 ? 64'hffffffffffffffff : 64'h0;
  assign T65 = T69 & T66;
  assign T66 = excSign ^ 1'h1;
  assign excSign = sign & T67;
  assign T67 = isNaN ^ 1'h1;
  assign isNaN = invalid & T68;
  assign T68 = exp[4'h9];
  assign T69 = io_signedOut ^ 1'h1;
  assign T70 = T74 | T77;
  assign T77 = {1'h0, T71};
  assign T71 = T72 ? 63'h7fffffffffffffff : 63'h0;
  assign T72 = io_signedOut & T73;
  assign T73 = excSign ^ 1'h1;
  assign T74 = T75 ? 64'h8000000000000000 : 64'h0;
  assign T75 = io_signedOut & excSign;
  assign T76 = invalid | overflow;
endmodule

module RecFNToIN_1(
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    input  io_signedOut,
    output[31:0] io_out,
    output[2:0] io_intExceptionFlags
);

  wire[2:0] T0;
  wire[1:0] T1;
  wire inexact;
  wire T2;
  wire T3;
  wire T4;
  wire roundInexact;
  wire T5;
  wire isZero;
  wire[2:0] T6;
  wire[11:0] exp;
  wire T7;
  wire[1:0] T8;
  wire[2:0] roundBits;
  wire T9;
  wire[50:0] T10;
  wire[83:0] shiftedSig;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[52:0] T13;
  wire[51:0] fract;
  wire[1:0] T14;
  wire notSpecial_magGeOne;
  wire overflow;
  wire overflow_unsigned;
  wire T15;
  wire roundIncr;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire roundIncr_nearestEven;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire T28;
  wire[10:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire sign;
  wire T36;
  wire T37;
  wire roundCarryBut2;
  wire T38;
  wire[29:0] T39;
  wire[31:0] unroundedInt;
  wire T40;
  wire T41;
  wire T42;
  wire[10:0] posExp;
  wire T43;
  wire T44;
  wire overflow_signed;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[30:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire invalid;
  wire[1:0] T59;
  wire[31:0] T60;
  wire[31:0] roundedInt;
  wire[31:0] complUnroundedInt;
  wire[31:0] T61;
  wire[31:0] T62;
  wire T63;
  wire[31:0] excValue;
  wire[31:0] T64;
  wire T65;
  wire T66;
  wire excSign;
  wire T67;
  wire isNaN;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire[31:0] T77;
  wire[30:0] T71;
  wire T72;
  wire T73;
  wire[31:0] T74;
  wire T75;
  wire T76;


  assign io_intExceptionFlags = T0;
  assign T0 = {invalid, T1};
  assign T1 = {overflow, inexact};
  assign inexact = T3 & T2;
  assign T2 = overflow ^ 1'h1;
  assign T3 = roundInexact & T4;
  assign T4 = invalid ^ 1'h1;
  assign roundInexact = notSpecial_magGeOne ? T7 : T5;
  assign T5 = isZero ^ 1'h1;
  assign isZero = T6 == 3'h0;
  assign T6 = exp[4'hb:4'h9];
  assign exp = io_in[6'h3f:6'h34];
  assign T7 = T8 != 2'h0;
  assign T8 = roundBits[1'h1:1'h0];
  assign roundBits = {T14, T9};
  assign T9 = T10 != 51'h0;
  assign T10 = shiftedSig[6'h32:1'h0];
  assign shiftedSig = T13 << T11;
  assign T11 = notSpecial_magGeOne ? T12 : 5'h0;
  assign T12 = exp[3'h4:1'h0];
  assign T13 = {notSpecial_magGeOne, fract};
  assign fract = io_in[6'h33:1'h0];
  assign T14 = shiftedSig[6'h34:6'h33];
  assign notSpecial_magGeOne = exp[4'hb];
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign overflow_unsigned = notSpecial_magGeOne ? T36 : T15;
  assign T15 = sign & roundIncr;
  assign roundIncr = T20 | T16;
  assign T16 = T19 & T17;
  assign T17 = T18 & roundInexact;
  assign T18 = sign ^ 1'h1;
  assign T19 = io_roundingMode == 2'h3;
  assign T20 = T24 | T21;
  assign T21 = T23 & T22;
  assign T22 = sign & roundInexact;
  assign T23 = io_roundingMode == 2'h2;
  assign T24 = T35 & roundIncr_nearestEven;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T30 : T25;
  assign T25 = T28 ? T26 : 1'h0;
  assign T26 = T27 != 2'h0;
  assign T27 = roundBits[1'h1:1'h0];
  assign T28 = T29 == 11'h7ff;
  assign T29 = exp[4'ha:1'h0];
  assign T30 = T33 | T31;
  assign T31 = T32 == 2'h3;
  assign T32 = roundBits[1'h1:1'h0];
  assign T33 = T34 == 2'h3;
  assign T34 = roundBits[2'h2:1'h1];
  assign T35 = io_roundingMode == 2'h0;
  assign sign = io_in[7'h40];
  assign T36 = T43 | T37;
  assign T37 = T40 & roundCarryBut2;
  assign roundCarryBut2 = T38 & roundIncr;
  assign T38 = T39 == 30'h3fffffff;
  assign T39 = unroundedInt[5'h1d:1'h0];
  assign unroundedInt = shiftedSig[7'h53:6'h34];
  assign T40 = T42 & T41;
  assign T41 = unroundedInt[5'h1e];
  assign T42 = posExp == 11'h1f;
  assign posExp = exp[4'ha:1'h0];
  assign T43 = sign | T44;
  assign T44 = 11'h20 <= posExp;
  assign overflow_signed = notSpecial_magGeOne ? T45 : 1'h0;
  assign T45 = T50 | T46;
  assign T46 = T47 & roundCarryBut2;
  assign T47 = T49 & T48;
  assign T48 = posExp == 11'h1e;
  assign T49 = sign ^ 1'h1;
  assign T50 = T58 | T51;
  assign T51 = T57 & T52;
  assign T52 = T53 | roundIncr;
  assign T53 = T56 | T54;
  assign T54 = T55 != 31'h0;
  assign T55 = unroundedInt[5'h1e:1'h0];
  assign T56 = sign ^ 1'h1;
  assign T57 = posExp == 11'h1f;
  assign T58 = 11'h20 <= posExp;
  assign invalid = T59 == 2'h3;
  assign T59 = exp[4'hb:4'ha];
  assign io_out = T60;
  assign T60 = T76 ? excValue : roundedInt;
  assign roundedInt = T63 ? T62 : complUnroundedInt;
  assign complUnroundedInt = sign ? T61 : unroundedInt;
  assign T61 = ~ unroundedInt;
  assign T62 = complUnroundedInt + 32'h1;
  assign T63 = roundIncr ^ sign;
  assign excValue = T70 | T64;
  assign T64 = T65 ? 32'hffffffff : 32'h0;
  assign T65 = T69 & T66;
  assign T66 = excSign ^ 1'h1;
  assign excSign = sign & T67;
  assign T67 = isNaN ^ 1'h1;
  assign isNaN = invalid & T68;
  assign T68 = exp[4'h9];
  assign T69 = io_signedOut ^ 1'h1;
  assign T70 = T74 | T77;
  assign T77 = {1'h0, T71};
  assign T71 = T72 ? 31'h7fffffff : 31'h0;
  assign T72 = io_signedOut & T73;
  assign T73 = excSign ^ 1'h1;
  assign T74 = T75 ? 32'h80000000 : 32'h0;
  assign T75 = io_signedOut & excSign;
  assign T76 = invalid | overflow;
endmodule

module FPToInt(input clk,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap12,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_div,
    input  io_in_bits_sqrt,
    input  io_in_bits_round,
    input  io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output[4:0] io_as_double_cmd,
    output io_as_double_ldst,
    output io_as_double_wen,
    output io_as_double_ren1,
    output io_as_double_ren2,
    output io_as_double_ren3,
    output io_as_double_swap12,
    output io_as_double_swap23,
    output io_as_double_single,
    output io_as_double_fromint,
    output io_as_double_toint,
    output io_as_double_fastpipe,
    output io_as_double_fma,
    output io_as_double_div,
    output io_as_double_sqrt,
    output io_as_double_round,
    output io_as_double_wflags,
    output[2:0] io_as_double_rm,
    output[1:0] io_as_double_typ,
    output[64:0] io_as_double_in1,
    output[64:0] io_as_double_in2,
    output[64:0] io_as_double_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output[63:0] io_out_bits_store,
    output[63:0] io_out_bits_toint,
    output[4:0] io_out_bits_exc
);

  wire T0;
  wire T1;
  reg [1:0] in_typ;
  wire[1:0] T2;
  wire[1:0] T227;
  reg [2:0] in_rm;
  wire[2:0] T3;
  reg [64:0] in_in1;
  wire[64:0] T4;
  wire[64:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] T228;
  reg [64:0] in_in2;
  wire[64:0] T15;
  wire[64:0] T16;
  wire[32:0] T229;
  wire[32:0] T230;
  wire[4:0] T17;
  wire[4:0] T18;
  wire T19;
  wire[4:0] T20;
  reg [4:0] in_cmd;
  wire[4:0] T21;
  wire[4:0] T22;
  wire[3:0] T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire T29;
  wire[4:0] T30;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[63:0] unrec_out;
  wire[63:0] unrec_d;
  wire[62:0] T34;
  wire[51:0] T35;
  wire[51:0] T36;
  wire[51:0] T37;
  wire[52:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[11:0] T41;
  wire[52:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[9:0] T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire[2:0] T50;
  wire[51:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  wire[10:0] T64;
  wire[10:0] T65;
  wire[10:0] T231;
  wire[10:0] T66;
  wire[10:0] T67;
  wire T68;
  wire[63:0] T69;
  wire[31:0] unrec_s;
  wire[30:0] T70;
  wire[22:0] T71;
  wire[22:0] T72;
  wire[22:0] T73;
  wire[23:0] T74;
  wire[4:0] T75;
  wire[4:0] T76;
  wire[8:0] T77;
  wire[23:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[6:0] T82;
  wire T83;
  wire[1:0] T84;
  wire T85;
  wire[2:0] T86;
  wire[22:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[1:0] T92;
  wire T93;
  wire T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire[1:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T232;
  wire[7:0] T102;
  wire[7:0] T103;
  wire T104;
  wire[31:0] T105;
  wire[31:0] T233;
  wire T106;
  reg  in_single;
  wire T107;
  wire[63:0] T234;
  wire[9:0] classify_out;
  wire[9:0] classify_d;
  wire[4:0] T108;
  wire[2:0] T109;
  wire[1:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[11:0] T116;
  wire T117;
  wire[1:0] T118;
  wire[2:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[9:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[1:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] T138;
  wire[2:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[51:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire[9:0] classify_s;
  wire[4:0] T155;
  wire[2:0] T156;
  wire[1:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[8:0] T163;
  wire T164;
  wire[1:0] T165;
  wire[2:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[6:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[4:0] T185;
  wire[2:0] T186;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire[22:0] T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[63:0] T235;
  wire dcmp_out;
  wire[2:0] T203;
  wire[2:0] T236;
  wire[1:0] T204;
  wire[2:0] T205;
  wire[63:0] T206;
  wire[63:0] T207;
  wire[63:0] T237;
  wire[31:0] T208;
  wire[31:0] T238;
  wire T239;
  wire[63:0] T209;
  wire T210;
  reg  valid;
  reg [64:0] in_in3;
  wire[64:0] T211;
  reg  in_wflags;
  wire T212;
  reg  in_round;
  wire T213;
  reg  in_sqrt;
  wire T214;
  reg  in_div;
  wire T215;
  reg  in_fma;
  wire T216;
  reg  in_fastpipe;
  wire T217;
  reg  in_toint;
  wire T218;
  reg  in_fromint;
  wire T219;
  reg  in_swap23;
  wire T220;
  reg  in_swap12;
  wire T221;
  reg  in_ren3;
  wire T222;
  reg  in_ren2;
  wire T223;
  reg  in_ren1;
  wire T224;
  reg  in_wen;
  wire T225;
  reg  in_ldst;
  wire T226;
  wire[64:0] RecFNToRecFN_io_out;
  wire[64:0] RecFNToRecFN_1_io_out;
  wire dcmp_io_lt;
  wire dcmp_io_eq;
  wire[4:0] dcmp_io_exceptionFlags;
  wire[63:0] d2l_io_out;
  wire[2:0] d2l_io_intExceptionFlags;
  wire[31:0] d2w_io_out;
  wire[2:0] d2w_io_intExceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_typ = {1{$random}};
    in_rm = {1{$random}};
    in_in1 = {3{$random}};
    in_in2 = {3{$random}};
    in_cmd = {1{$random}};
    in_single = {1{$random}};
    valid = {1{$random}};
    in_in3 = {3{$random}};
    in_wflags = {1{$random}};
    in_round = {1{$random}};
    in_sqrt = {1{$random}};
    in_div = {1{$random}};
    in_fma = {1{$random}};
    in_fastpipe = {1{$random}};
    in_toint = {1{$random}};
    in_fromint = {1{$random}};
    in_swap23 = {1{$random}};
    in_swap12 = {1{$random}};
    in_ren3 = {1{$random}};
    in_ren2 = {1{$random}};
    in_ren1 = {1{$random}};
    in_wen = {1{$random}};
    in_ldst = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = ~ T1;
  assign T1 = in_typ[1'h0];
  assign T2 = io_in_valid ? io_in_bits_typ : in_typ;
  assign T227 = in_rm[1'h1:1'h0];
  assign T3 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T4 = T6 ? RecFNToRecFN_io_out : T5;
  assign T5 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T6 = io_in_valid & T7;
  assign T7 = T11 & T8;
  assign T8 = T9 ^ 1'h1;
  assign T9 = 5'hc == T10;
  assign T10 = io_in_bits_cmd & 5'hc;
  assign T11 = io_in_bits_single & T12;
  assign T12 = io_in_bits_ldst ^ 1'h1;
  assign T13 = ~ T14;
  assign T14 = in_typ[1'h0];
  assign T228 = in_rm[1'h1:1'h0];
  assign T15 = T6 ? RecFNToRecFN_1_io_out : T16;
  assign T16 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T229 = io_in_bits_in2[6'h20:1'h0];
  assign T230 = io_in_bits_in1[6'h20:1'h0];
  assign io_out_bits_exc = T17;
  assign T17 = T29 ? T22 : T18;
  assign T18 = T19 ? dcmp_io_exceptionFlags : 5'h0;
  assign T19 = 5'h4 == T20;
  assign T20 = in_cmd & 5'hc;
  assign T21 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T22 = {T27, T23};
  assign T23 = {3'h0, T24};
  assign T24 = T25[1'h0];
  assign T25 = T26 ? d2l_io_intExceptionFlags : d2w_io_intExceptionFlags;
  assign T26 = in_typ[1'h1];
  assign T27 = T28 != 2'h0;
  assign T28 = T25[2'h2:1'h1];
  assign T29 = 5'h8 == T30;
  assign T30 = in_cmd & 5'hc;
  assign io_out_bits_toint = T31;
  assign T31 = T29 ? T206 : T32;
  assign T32 = T19 ? T235 : T33;
  assign T33 = T202 ? T234 : unrec_out;
  assign unrec_out = in_single ? T69 : unrec_d;
  assign unrec_d = {T68, T34};
  assign T34 = {T64, T35};
  assign T35 = T52 ? T51 : T36;
  assign T36 = T43 ? T37 : 52'h0;
  assign T37 = T38[6'h33:1'h0];
  assign T38 = T42 >> T39;
  assign T39 = 6'h2 - T40;
  assign T40 = T41[3'h5:1'h0];
  assign T41 = in_in1[6'h3f:6'h34];
  assign T42 = {1'h1, T51};
  assign T43 = T49 | T44;
  assign T44 = T47 & T45;
  assign T45 = T46 < 10'h2;
  assign T46 = T41[4'h9:1'h0];
  assign T47 = T48 == 2'h1;
  assign T48 = T41[4'hb:4'ha];
  assign T49 = T50 == 3'h1;
  assign T50 = T41[4'hb:4'h9];
  assign T51 = in_in1[6'h33:1'h0];
  assign T52 = T57 | T53;
  assign T53 = T55 & T54;
  assign T54 = T41[4'h9];
  assign T55 = T56 == 2'h3;
  assign T56 = T41[4'hb:4'ha];
  assign T57 = T60 | T58;
  assign T58 = T59 == 2'h2;
  assign T59 = T41[4'hb:4'ha];
  assign T60 = T62 & T61;
  assign T61 = T45 ^ 1'h1;
  assign T62 = T63 == 2'h1;
  assign T63 = T41[4'hb:4'ha];
  assign T64 = T57 ? T66 : T65;
  assign T65 = 11'h0 - T231;
  assign T231 = {10'h0, T55};
  assign T66 = T67 - 11'h401;
  assign T67 = T41[4'ha:1'h0];
  assign T68 = in_in1[7'h40];
  assign T69 = {T105, unrec_s};
  assign unrec_s = {T104, T70};
  assign T70 = {T100, T71};
  assign T71 = T88 ? T87 : T72;
  assign T72 = T79 ? T73 : 23'h0;
  assign T73 = T74[5'h16:1'h0];
  assign T74 = T78 >> T75;
  assign T75 = 5'h2 - T76;
  assign T76 = T77[3'h4:1'h0];
  assign T77 = in_in1[5'h1f:5'h17];
  assign T78 = {1'h1, T87};
  assign T79 = T85 | T80;
  assign T80 = T83 & T81;
  assign T81 = T82 < 7'h2;
  assign T82 = T77[3'h6:1'h0];
  assign T83 = T84 == 2'h1;
  assign T84 = T77[4'h8:3'h7];
  assign T85 = T86 == 3'h1;
  assign T86 = T77[4'h8:3'h6];
  assign T87 = in_in1[5'h16:1'h0];
  assign T88 = T93 | T89;
  assign T89 = T91 & T90;
  assign T90 = T77[3'h6];
  assign T91 = T92 == 2'h3;
  assign T92 = T77[4'h8:3'h7];
  assign T93 = T96 | T94;
  assign T94 = T95 == 2'h2;
  assign T95 = T77[4'h8:3'h7];
  assign T96 = T98 & T97;
  assign T97 = T81 ^ 1'h1;
  assign T98 = T99 == 2'h1;
  assign T99 = T77[4'h8:3'h7];
  assign T100 = T93 ? T102 : T101;
  assign T101 = 8'h0 - T232;
  assign T232 = {7'h0, T91};
  assign T102 = T103 - 8'h81;
  assign T103 = T77[3'h7:1'h0];
  assign T104 = in_in1[6'h20];
  assign T105 = 32'h0 - T233;
  assign T233 = {31'h0, T106};
  assign T106 = unrec_s[5'h1f];
  assign T107 = io_in_valid ? io_in_bits_single : in_single;
  assign T234 = {54'h0, classify_out};
  assign classify_out = in_single ? classify_s : classify_d;
  assign classify_d = {T138, T108};
  assign T108 = {T133, T109};
  assign T109 = {T128, T110};
  assign T110 = {T120, T111};
  assign T111 = T113 & T112;
  assign T112 = in_in1[7'h40];
  assign T113 = T117 & T114;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116[4'h9];
  assign T116 = in_in1[6'h3f:6'h34];
  assign T117 = T118 == 2'h3;
  assign T118 = T119[2'h2:1'h1];
  assign T119 = T116[4'hb:4'h9];
  assign T120 = T121 & T112;
  assign T121 = T123 | T122;
  assign T122 = T118 == 2'h2;
  assign T123 = T127 & T124;
  assign T124 = T125 ^ 1'h1;
  assign T125 = T126 < 10'h2;
  assign T126 = T116[4'h9:1'h0];
  assign T127 = T118 == 2'h1;
  assign T128 = T129 & T112;
  assign T129 = T132 | T130;
  assign T130 = T131 & T125;
  assign T131 = T118 == 2'h1;
  assign T132 = T119 == 3'h1;
  assign T133 = {T136, T134};
  assign T134 = T135 & T112;
  assign T135 = T119 == 3'h0;
  assign T136 = T135 & T137;
  assign T137 = T112 ^ 1'h1;
  assign T138 = {T147, T139};
  assign T139 = {T145, T140};
  assign T140 = {T143, T141};
  assign T141 = T129 & T142;
  assign T142 = T112 ^ 1'h1;
  assign T143 = T121 & T144;
  assign T144 = T112 ^ 1'h1;
  assign T145 = T113 & T146;
  assign T146 = T112 ^ 1'h1;
  assign T147 = {T153, T148};
  assign T148 = T152 & T149;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T151[6'h33];
  assign T151 = in_in1[6'h33:1'h0];
  assign T152 = T119 == 3'h7;
  assign T153 = T152 & T154;
  assign T154 = T151[6'h33];
  assign classify_s = {T185, T155};
  assign T155 = {T180, T156};
  assign T156 = {T175, T157};
  assign T157 = {T167, T158};
  assign T158 = T160 & T159;
  assign T159 = in_in1[6'h20];
  assign T160 = T164 & T161;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T163[3'h6];
  assign T163 = in_in1[5'h1f:5'h17];
  assign T164 = T165 == 2'h3;
  assign T165 = T166[2'h2:1'h1];
  assign T166 = T163[4'h8:3'h6];
  assign T167 = T168 & T159;
  assign T168 = T170 | T169;
  assign T169 = T165 == 2'h2;
  assign T170 = T174 & T171;
  assign T171 = T172 ^ 1'h1;
  assign T172 = T173 < 7'h2;
  assign T173 = T163[3'h6:1'h0];
  assign T174 = T165 == 2'h1;
  assign T175 = T176 & T159;
  assign T176 = T179 | T177;
  assign T177 = T178 & T172;
  assign T178 = T165 == 2'h1;
  assign T179 = T166 == 3'h1;
  assign T180 = {T183, T181};
  assign T181 = T182 & T159;
  assign T182 = T166 == 3'h0;
  assign T183 = T182 & T184;
  assign T184 = T159 ^ 1'h1;
  assign T185 = {T194, T186};
  assign T186 = {T192, T187};
  assign T187 = {T190, T188};
  assign T188 = T176 & T189;
  assign T189 = T159 ^ 1'h1;
  assign T190 = T168 & T191;
  assign T191 = T159 ^ 1'h1;
  assign T192 = T160 & T193;
  assign T193 = T159 ^ 1'h1;
  assign T194 = {T200, T195};
  assign T195 = T199 & T196;
  assign T196 = T197 ^ 1'h1;
  assign T197 = T198[5'h16];
  assign T198 = in_in1[5'h16:1'h0];
  assign T199 = T166 == 3'h7;
  assign T200 = T199 & T201;
  assign T201 = T198[5'h16];
  assign T202 = in_rm[1'h0];
  assign T235 = {63'h0, dcmp_out};
  assign dcmp_out = T203 != 3'h0;
  assign T203 = T205 & T236;
  assign T236 = {1'h0, T204};
  assign T204 = {dcmp_io_lt, dcmp_io_eq};
  assign T205 = ~ in_rm;
  assign T206 = T207;
  assign T207 = T210 ? T209 : T237;
  assign T237 = {T238, T208};
  assign T208 = d2w_io_out;
  assign T238 = T239 ? 32'hffffffff : 32'h0;
  assign T239 = T208[5'h1f];
  assign T209 = d2l_io_out;
  assign T210 = in_typ[1'h1];
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_lt = dcmp_io_lt;
  assign io_out_valid = valid;
  assign io_as_double_in3 = in_in3;
  assign T211 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign io_as_double_in2 = in_in2;
  assign io_as_double_in1 = in_in1;
  assign io_as_double_typ = in_typ;
  assign io_as_double_rm = in_rm;
  assign io_as_double_wflags = in_wflags;
  assign T212 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign io_as_double_round = in_round;
  assign T213 = io_in_valid ? io_in_bits_round : in_round;
  assign io_as_double_sqrt = in_sqrt;
  assign T214 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign io_as_double_div = in_div;
  assign T215 = io_in_valid ? io_in_bits_div : in_div;
  assign io_as_double_fma = in_fma;
  assign T216 = io_in_valid ? io_in_bits_fma : in_fma;
  assign io_as_double_fastpipe = in_fastpipe;
  assign T217 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign io_as_double_toint = in_toint;
  assign T218 = io_in_valid ? io_in_bits_toint : in_toint;
  assign io_as_double_fromint = in_fromint;
  assign T219 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign io_as_double_single = in_single;
  assign io_as_double_swap23 = in_swap23;
  assign T220 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign io_as_double_swap12 = in_swap12;
  assign T221 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign io_as_double_ren3 = in_ren3;
  assign T222 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign io_as_double_ren2 = in_ren2;
  assign T223 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign io_as_double_ren1 = in_ren1;
  assign T224 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign io_as_double_wen = in_wen;
  assign T225 = io_in_valid ? io_in_bits_wen : in_wen;
  assign io_as_double_ldst = in_ldst;
  assign T226 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign io_as_double_cmd = in_cmd;
  RecFNToRecFN RecFNToRecFN(
       .io_in( T230 ),
       .io_roundingMode( 2'h0 ),
       .io_out( RecFNToRecFN_io_out )
       //.io_exceptionFlags(  )
  );
  RecFNToRecFN RecFNToRecFN_1(
       .io_in( T229 ),
       .io_roundingMode( 2'h0 ),
       .io_out( RecFNToRecFN_1_io_out )
       //.io_exceptionFlags(  )
  );
  CompareRecFN dcmp(
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_signaling( 1'h1 ),
       .io_lt( dcmp_io_lt ),
       .io_eq( dcmp_io_eq ),
       //.io_gt(  )
       .io_exceptionFlags( dcmp_io_exceptionFlags )
  );
  RecFNToIN_0 d2l(
       .io_in( in_in1 ),
       .io_roundingMode( T228 ),
       .io_signedOut( T13 ),
       .io_out( d2l_io_out ),
       .io_intExceptionFlags( d2l_io_intExceptionFlags )
  );
  RecFNToIN_1 d2w(
       .io_in( in_in1 ),
       .io_roundingMode( T227 ),
       .io_signedOut( T0 ),
       .io_out( d2w_io_out ),
       .io_intExceptionFlags( d2w_io_intExceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T6) begin
      in_in1 <= RecFNToRecFN_io_out;
    end else if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(T6) begin
      in_in2 <= RecFNToRecFN_1_io_out;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      in_single <= io_in_bits_single;
    end
    valid <= io_in_valid;
    if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(io_in_valid) begin
      in_wflags <= io_in_bits_wflags;
    end
    if(io_in_valid) begin
      in_round <= io_in_bits_round;
    end
    if(io_in_valid) begin
      in_sqrt <= io_in_bits_sqrt;
    end
    if(io_in_valid) begin
      in_div <= io_in_bits_div;
    end
    if(io_in_valid) begin
      in_fma <= io_in_bits_fma;
    end
    if(io_in_valid) begin
      in_fastpipe <= io_in_bits_fastpipe;
    end
    if(io_in_valid) begin
      in_toint <= io_in_bits_toint;
    end
    if(io_in_valid) begin
      in_fromint <= io_in_bits_fromint;
    end
    if(io_in_valid) begin
      in_swap23 <= io_in_bits_swap23;
    end
    if(io_in_valid) begin
      in_swap12 <= io_in_bits_swap12;
    end
    if(io_in_valid) begin
      in_ren3 <= io_in_bits_ren3;
    end
    if(io_in_valid) begin
      in_ren2 <= io_in_bits_ren2;
    end
    if(io_in_valid) begin
      in_ren1 <= io_in_bits_ren1;
    end
    if(io_in_valid) begin
      in_wen <= io_in_bits_wen;
    end
    if(io_in_valid) begin
      in_ldst <= io_in_bits_ldst;
    end
  end
endmodule

module INToRecFN_0(
    input  io_signedIn,
    input [63:0] io_in,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[1:0] T1;
  wire inexact;
  wire[1:0] T2;
  wire[2:0] roundBits;
  wire T3;
  wire[38:0] T4;
  wire[63:0] normAbsIn;
  wire[126:0] T5;
  wire[5:0] normCount;
  wire[5:0] T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire[5:0] T48;
  wire[5:0] T49;
  wire[5:0] T50;
  wire[5:0] T51;
  wire[5:0] T52;
  wire[5:0] T53;
  wire[5:0] T54;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire[5:0] T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[4:0] T69;
  wire[4:0] T70;
  wire[4:0] T71;
  wire[4:0] T72;
  wire[4:0] T73;
  wire[4:0] T74;
  wire[4:0] T75;
  wire[4:0] T76;
  wire[4:0] T77;
  wire[4:0] T78;
  wire[4:0] T79;
  wire[4:0] T80;
  wire[4:0] T81;
  wire[4:0] T82;
  wire[4:0] T83;
  wire[4:0] T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire[3:0] T87;
  wire[3:0] T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire[63:0] T7;
  wire[63:0] T8;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[63:0] absIn;
  wire[63:0] T9;
  wire sign;
  wire T10;
  wire[1:0] T11;
  wire[32:0] T12;
  wire[31:0] T13;
  wire[22:0] T14;
  wire[24:0] roundedNorm;
  wire[24:0] unroundedNorm;
  wire[23:0] T15;
  wire[24:0] T16;
  wire round;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire T29;
  wire[1:0] T30;
  wire T31;
  wire[8:0] expOut;
  wire[7:0] T32;
  wire[7:0] roundedExp;
  wire[7:0] T162;
  wire T33;
  wire[7:0] T34;
  wire[6:0] unroundedExp;
  wire[5:0] T35;
  wire T36;


  assign io_exceptionFlags = T0;
  assign T0 = {3'h0, T1};
  assign T1 = {1'h0, inexact};
  assign inexact = T2 != 2'h0;
  assign T2 = roundBits[1'h1:1'h0];
  assign roundBits = {T11, T3};
  assign T3 = T4 != 39'h0;
  assign T4 = normAbsIn[6'h26:1'h0];
  assign normAbsIn = T5[6'h3f:1'h0];
  assign T5 = absIn << normCount;
  assign normCount = ~ T37;
  assign T37 = T161 ? 6'h3f : T38;
  assign T38 = T160 ? 6'h3e : T39;
  assign T39 = T159 ? 6'h3d : T40;
  assign T40 = T158 ? 6'h3c : T41;
  assign T41 = T157 ? 6'h3b : T42;
  assign T42 = T156 ? 6'h3a : T43;
  assign T43 = T155 ? 6'h39 : T44;
  assign T44 = T154 ? 6'h38 : T45;
  assign T45 = T153 ? 6'h37 : T46;
  assign T46 = T152 ? 6'h36 : T47;
  assign T47 = T151 ? 6'h35 : T48;
  assign T48 = T150 ? 6'h34 : T49;
  assign T49 = T149 ? 6'h33 : T50;
  assign T50 = T148 ? 6'h32 : T51;
  assign T51 = T147 ? 6'h31 : T52;
  assign T52 = T146 ? 6'h30 : T53;
  assign T53 = T145 ? 6'h2f : T54;
  assign T54 = T144 ? 6'h2e : T55;
  assign T55 = T143 ? 6'h2d : T56;
  assign T56 = T142 ? 6'h2c : T57;
  assign T57 = T141 ? 6'h2b : T58;
  assign T58 = T140 ? 6'h2a : T59;
  assign T59 = T139 ? 6'h29 : T60;
  assign T60 = T138 ? 6'h28 : T61;
  assign T61 = T137 ? 6'h27 : T62;
  assign T62 = T136 ? 6'h26 : T63;
  assign T63 = T135 ? 6'h25 : T64;
  assign T64 = T134 ? 6'h24 : T65;
  assign T65 = T133 ? 6'h23 : T66;
  assign T66 = T132 ? 6'h22 : T67;
  assign T67 = T131 ? 6'h21 : T68;
  assign T68 = T130 ? 6'h20 : T69;
  assign T69 = T129 ? 5'h1f : T70;
  assign T70 = T128 ? 5'h1e : T71;
  assign T71 = T127 ? 5'h1d : T72;
  assign T72 = T126 ? 5'h1c : T73;
  assign T73 = T125 ? 5'h1b : T74;
  assign T74 = T124 ? 5'h1a : T75;
  assign T75 = T123 ? 5'h19 : T76;
  assign T76 = T122 ? 5'h18 : T77;
  assign T77 = T121 ? 5'h17 : T78;
  assign T78 = T120 ? 5'h16 : T79;
  assign T79 = T119 ? 5'h15 : T80;
  assign T80 = T118 ? 5'h14 : T81;
  assign T81 = T117 ? 5'h13 : T82;
  assign T82 = T116 ? 5'h12 : T83;
  assign T83 = T115 ? 5'h11 : T84;
  assign T84 = T114 ? 5'h10 : T85;
  assign T85 = T113 ? 4'hf : T86;
  assign T86 = T112 ? 4'he : T87;
  assign T87 = T111 ? 4'hd : T88;
  assign T88 = T110 ? 4'hc : T89;
  assign T89 = T109 ? 4'hb : T90;
  assign T90 = T108 ? 4'ha : T91;
  assign T91 = T107 ? 4'h9 : T92;
  assign T92 = T106 ? 4'h8 : T93;
  assign T93 = T105 ? 3'h7 : T94;
  assign T94 = T104 ? 3'h6 : T95;
  assign T95 = T103 ? 3'h5 : T96;
  assign T96 = T102 ? 3'h4 : T97;
  assign T97 = T101 ? 2'h3 : T98;
  assign T98 = T100 ? 2'h2 : T99;
  assign T99 = T7[1'h1];
  assign T7 = T8;
  assign T8 = absIn << 1'h0;
  assign T100 = T7[2'h2];
  assign T101 = T7[2'h3];
  assign T102 = T7[3'h4];
  assign T103 = T7[3'h5];
  assign T104 = T7[3'h6];
  assign T105 = T7[3'h7];
  assign T106 = T7[4'h8];
  assign T107 = T7[4'h9];
  assign T108 = T7[4'ha];
  assign T109 = T7[4'hb];
  assign T110 = T7[4'hc];
  assign T111 = T7[4'hd];
  assign T112 = T7[4'he];
  assign T113 = T7[4'hf];
  assign T114 = T7[5'h10];
  assign T115 = T7[5'h11];
  assign T116 = T7[5'h12];
  assign T117 = T7[5'h13];
  assign T118 = T7[5'h14];
  assign T119 = T7[5'h15];
  assign T120 = T7[5'h16];
  assign T121 = T7[5'h17];
  assign T122 = T7[5'h18];
  assign T123 = T7[5'h19];
  assign T124 = T7[5'h1a];
  assign T125 = T7[5'h1b];
  assign T126 = T7[5'h1c];
  assign T127 = T7[5'h1d];
  assign T128 = T7[5'h1e];
  assign T129 = T7[5'h1f];
  assign T130 = T7[6'h20];
  assign T131 = T7[6'h21];
  assign T132 = T7[6'h22];
  assign T133 = T7[6'h23];
  assign T134 = T7[6'h24];
  assign T135 = T7[6'h25];
  assign T136 = T7[6'h26];
  assign T137 = T7[6'h27];
  assign T138 = T7[6'h28];
  assign T139 = T7[6'h29];
  assign T140 = T7[6'h2a];
  assign T141 = T7[6'h2b];
  assign T142 = T7[6'h2c];
  assign T143 = T7[6'h2d];
  assign T144 = T7[6'h2e];
  assign T145 = T7[6'h2f];
  assign T146 = T7[6'h30];
  assign T147 = T7[6'h31];
  assign T148 = T7[6'h32];
  assign T149 = T7[6'h33];
  assign T150 = T7[6'h34];
  assign T151 = T7[6'h35];
  assign T152 = T7[6'h36];
  assign T153 = T7[6'h37];
  assign T154 = T7[6'h38];
  assign T155 = T7[6'h39];
  assign T156 = T7[6'h3a];
  assign T157 = T7[6'h3b];
  assign T158 = T7[6'h3c];
  assign T159 = T7[6'h3d];
  assign T160 = T7[6'h3e];
  assign T161 = T7[6'h3f];
  assign absIn = sign ? T9 : io_in;
  assign T9 = 64'h0 - io_in;
  assign sign = io_signedIn & T10;
  assign T10 = io_in[6'h3f];
  assign T11 = normAbsIn[6'h28:6'h27];
  assign io_out = T12;
  assign T12 = {sign, T13};
  assign T13 = {expOut, T14};
  assign T14 = roundedNorm[5'h16:1'h0];
  assign roundedNorm = round ? T16 : unroundedNorm;
  assign unroundedNorm = {1'h0, T15};
  assign T15 = normAbsIn[6'h3f:6'h28];
  assign T16 = unroundedNorm + 25'h1;
  assign round = T21 | T17;
  assign T17 = T20 ? T18 : 1'h0;
  assign T18 = T19 & inexact;
  assign T19 = sign ^ 1'h1;
  assign T20 = io_roundingMode == 2'h3;
  assign T21 = T25 | T22;
  assign T22 = T24 ? T23 : 1'h0;
  assign T23 = sign & inexact;
  assign T24 = io_roundingMode == 2'h2;
  assign T25 = T31 ? T26 : 1'h0;
  assign T26 = T29 | T27;
  assign T27 = T28 == 2'h3;
  assign T28 = roundBits[1'h1:1'h0];
  assign T29 = T30 == 2'h3;
  assign T30 = roundBits[2'h2:1'h1];
  assign T31 = io_roundingMode == 2'h0;
  assign expOut = {T36, T32};
  assign T32 = roundedExp;
  assign roundedExp = T34 + T162;
  assign T162 = {7'h0, T33};
  assign T33 = roundedNorm[5'h18];
  assign T34 = {1'h0, unroundedExp};
  assign unroundedExp = {1'h0, T35};
  assign T35 = ~ normCount;
  assign T36 = normAbsIn[6'h3f];
endmodule

module INToRecFN_1(
    input  io_signedIn,
    input [63:0] io_in,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[1:0] T1;
  wire inexact;
  wire[1:0] T2;
  wire[2:0] roundBits;
  wire T3;
  wire[9:0] T4;
  wire[63:0] normAbsIn;
  wire[126:0] T5;
  wire[5:0] normCount;
  wire[5:0] T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire[5:0] T48;
  wire[5:0] T49;
  wire[5:0] T50;
  wire[5:0] T51;
  wire[5:0] T52;
  wire[5:0] T53;
  wire[5:0] T54;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire[5:0] T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[4:0] T69;
  wire[4:0] T70;
  wire[4:0] T71;
  wire[4:0] T72;
  wire[4:0] T73;
  wire[4:0] T74;
  wire[4:0] T75;
  wire[4:0] T76;
  wire[4:0] T77;
  wire[4:0] T78;
  wire[4:0] T79;
  wire[4:0] T80;
  wire[4:0] T81;
  wire[4:0] T82;
  wire[4:0] T83;
  wire[4:0] T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire[3:0] T87;
  wire[3:0] T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire[2:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire[63:0] T7;
  wire[63:0] T8;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[63:0] absIn;
  wire[63:0] T9;
  wire sign;
  wire T10;
  wire[1:0] T11;
  wire[64:0] T12;
  wire[63:0] T13;
  wire[51:0] T14;
  wire[53:0] roundedNorm;
  wire[53:0] unroundedNorm;
  wire[52:0] T15;
  wire[53:0] T16;
  wire round;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire T29;
  wire[1:0] T30;
  wire T31;
  wire[11:0] expOut;
  wire[10:0] T32;
  wire[10:0] roundedExp;
  wire[10:0] T162;
  wire T33;
  wire[10:0] T34;
  wire[9:0] unroundedExp;
  wire[5:0] T35;
  wire T36;


  assign io_exceptionFlags = T0;
  assign T0 = {3'h0, T1};
  assign T1 = {1'h0, inexact};
  assign inexact = T2 != 2'h0;
  assign T2 = roundBits[1'h1:1'h0];
  assign roundBits = {T11, T3};
  assign T3 = T4 != 10'h0;
  assign T4 = normAbsIn[4'h9:1'h0];
  assign normAbsIn = T5[6'h3f:1'h0];
  assign T5 = absIn << normCount;
  assign normCount = ~ T37;
  assign T37 = T161 ? 6'h3f : T38;
  assign T38 = T160 ? 6'h3e : T39;
  assign T39 = T159 ? 6'h3d : T40;
  assign T40 = T158 ? 6'h3c : T41;
  assign T41 = T157 ? 6'h3b : T42;
  assign T42 = T156 ? 6'h3a : T43;
  assign T43 = T155 ? 6'h39 : T44;
  assign T44 = T154 ? 6'h38 : T45;
  assign T45 = T153 ? 6'h37 : T46;
  assign T46 = T152 ? 6'h36 : T47;
  assign T47 = T151 ? 6'h35 : T48;
  assign T48 = T150 ? 6'h34 : T49;
  assign T49 = T149 ? 6'h33 : T50;
  assign T50 = T148 ? 6'h32 : T51;
  assign T51 = T147 ? 6'h31 : T52;
  assign T52 = T146 ? 6'h30 : T53;
  assign T53 = T145 ? 6'h2f : T54;
  assign T54 = T144 ? 6'h2e : T55;
  assign T55 = T143 ? 6'h2d : T56;
  assign T56 = T142 ? 6'h2c : T57;
  assign T57 = T141 ? 6'h2b : T58;
  assign T58 = T140 ? 6'h2a : T59;
  assign T59 = T139 ? 6'h29 : T60;
  assign T60 = T138 ? 6'h28 : T61;
  assign T61 = T137 ? 6'h27 : T62;
  assign T62 = T136 ? 6'h26 : T63;
  assign T63 = T135 ? 6'h25 : T64;
  assign T64 = T134 ? 6'h24 : T65;
  assign T65 = T133 ? 6'h23 : T66;
  assign T66 = T132 ? 6'h22 : T67;
  assign T67 = T131 ? 6'h21 : T68;
  assign T68 = T130 ? 6'h20 : T69;
  assign T69 = T129 ? 5'h1f : T70;
  assign T70 = T128 ? 5'h1e : T71;
  assign T71 = T127 ? 5'h1d : T72;
  assign T72 = T126 ? 5'h1c : T73;
  assign T73 = T125 ? 5'h1b : T74;
  assign T74 = T124 ? 5'h1a : T75;
  assign T75 = T123 ? 5'h19 : T76;
  assign T76 = T122 ? 5'h18 : T77;
  assign T77 = T121 ? 5'h17 : T78;
  assign T78 = T120 ? 5'h16 : T79;
  assign T79 = T119 ? 5'h15 : T80;
  assign T80 = T118 ? 5'h14 : T81;
  assign T81 = T117 ? 5'h13 : T82;
  assign T82 = T116 ? 5'h12 : T83;
  assign T83 = T115 ? 5'h11 : T84;
  assign T84 = T114 ? 5'h10 : T85;
  assign T85 = T113 ? 4'hf : T86;
  assign T86 = T112 ? 4'he : T87;
  assign T87 = T111 ? 4'hd : T88;
  assign T88 = T110 ? 4'hc : T89;
  assign T89 = T109 ? 4'hb : T90;
  assign T90 = T108 ? 4'ha : T91;
  assign T91 = T107 ? 4'h9 : T92;
  assign T92 = T106 ? 4'h8 : T93;
  assign T93 = T105 ? 3'h7 : T94;
  assign T94 = T104 ? 3'h6 : T95;
  assign T95 = T103 ? 3'h5 : T96;
  assign T96 = T102 ? 3'h4 : T97;
  assign T97 = T101 ? 2'h3 : T98;
  assign T98 = T100 ? 2'h2 : T99;
  assign T99 = T7[1'h1];
  assign T7 = T8;
  assign T8 = absIn << 1'h0;
  assign T100 = T7[2'h2];
  assign T101 = T7[2'h3];
  assign T102 = T7[3'h4];
  assign T103 = T7[3'h5];
  assign T104 = T7[3'h6];
  assign T105 = T7[3'h7];
  assign T106 = T7[4'h8];
  assign T107 = T7[4'h9];
  assign T108 = T7[4'ha];
  assign T109 = T7[4'hb];
  assign T110 = T7[4'hc];
  assign T111 = T7[4'hd];
  assign T112 = T7[4'he];
  assign T113 = T7[4'hf];
  assign T114 = T7[5'h10];
  assign T115 = T7[5'h11];
  assign T116 = T7[5'h12];
  assign T117 = T7[5'h13];
  assign T118 = T7[5'h14];
  assign T119 = T7[5'h15];
  assign T120 = T7[5'h16];
  assign T121 = T7[5'h17];
  assign T122 = T7[5'h18];
  assign T123 = T7[5'h19];
  assign T124 = T7[5'h1a];
  assign T125 = T7[5'h1b];
  assign T126 = T7[5'h1c];
  assign T127 = T7[5'h1d];
  assign T128 = T7[5'h1e];
  assign T129 = T7[5'h1f];
  assign T130 = T7[6'h20];
  assign T131 = T7[6'h21];
  assign T132 = T7[6'h22];
  assign T133 = T7[6'h23];
  assign T134 = T7[6'h24];
  assign T135 = T7[6'h25];
  assign T136 = T7[6'h26];
  assign T137 = T7[6'h27];
  assign T138 = T7[6'h28];
  assign T139 = T7[6'h29];
  assign T140 = T7[6'h2a];
  assign T141 = T7[6'h2b];
  assign T142 = T7[6'h2c];
  assign T143 = T7[6'h2d];
  assign T144 = T7[6'h2e];
  assign T145 = T7[6'h2f];
  assign T146 = T7[6'h30];
  assign T147 = T7[6'h31];
  assign T148 = T7[6'h32];
  assign T149 = T7[6'h33];
  assign T150 = T7[6'h34];
  assign T151 = T7[6'h35];
  assign T152 = T7[6'h36];
  assign T153 = T7[6'h37];
  assign T154 = T7[6'h38];
  assign T155 = T7[6'h39];
  assign T156 = T7[6'h3a];
  assign T157 = T7[6'h3b];
  assign T158 = T7[6'h3c];
  assign T159 = T7[6'h3d];
  assign T160 = T7[6'h3e];
  assign T161 = T7[6'h3f];
  assign absIn = sign ? T9 : io_in;
  assign T9 = 64'h0 - io_in;
  assign sign = io_signedIn & T10;
  assign T10 = io_in[6'h3f];
  assign T11 = normAbsIn[4'hb:4'ha];
  assign io_out = T12;
  assign T12 = {sign, T13};
  assign T13 = {expOut, T14};
  assign T14 = roundedNorm[6'h33:1'h0];
  assign roundedNorm = round ? T16 : unroundedNorm;
  assign unroundedNorm = {1'h0, T15};
  assign T15 = normAbsIn[6'h3f:4'hb];
  assign T16 = unroundedNorm + 54'h1;
  assign round = T21 | T17;
  assign T17 = T20 ? T18 : 1'h0;
  assign T18 = T19 & inexact;
  assign T19 = sign ^ 1'h1;
  assign T20 = io_roundingMode == 2'h3;
  assign T21 = T25 | T22;
  assign T22 = T24 ? T23 : 1'h0;
  assign T23 = sign & inexact;
  assign T24 = io_roundingMode == 2'h2;
  assign T25 = T31 ? T26 : 1'h0;
  assign T26 = T29 | T27;
  assign T27 = T28 == 2'h3;
  assign T28 = roundBits[1'h1:1'h0];
  assign T29 = T30 == 2'h3;
  assign T30 = roundBits[2'h2:1'h1];
  assign T31 = io_roundingMode == 2'h0;
  assign expOut = {T36, T32};
  assign T32 = roundedExp;
  assign roundedExp = T34 + T162;
  assign T162 = {10'h0, T33};
  assign T33 = roundedNorm[6'h35];
  assign T34 = {1'h0, unroundedExp};
  assign unroundedExp = {4'h0, T35};
  assign T35 = ~ normCount;
  assign T36 = normAbsIn[6'h3f];
endmodule

module IntToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap12,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_div,
    input  io_in_bits_sqrt,
    input  io_in_bits_round,
    input  io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T110;
  reg [2:0] R0;
  wire[2:0] T1;
  wire[63:0] T111;
  wire[64:0] T2;
  wire[64:0] longValue;
  wire[64:0] T112;
  wire[32:0] T3;
  wire[32:0] T113;
  wire[31:0] T4;
  wire[31:0] T5;
  reg [64:0] R6;
  wire[64:0] T7;
  wire T114;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[31:0] T10;
  wire T11;
  reg [1:0] R12;
  wire[1:0] T13;
  wire[31:0] T115;
  wire T116;
  wire[64:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire[1:0] T117;
  wire[63:0] T118;
  wire[64:0] T18;
  wire T19;
  wire T20;
  reg [4:0] R21;
  wire[4:0] T22;
  reg [4:0] R23;
  wire[4:0] T24;
  wire[4:0] mux_exc;
  wire[4:0] T25;
  wire[4:0] T26;
  wire T27;
  reg  R28;
  wire T29;
  wire T30;
  wire[4:0] T31;
  reg [4:0] R32;
  wire[4:0] T33;
  wire T34;
  wire T35;
  reg  R36;
  wire T119;
  reg  R37;
  wire T120;
  reg [64:0] R38;
  wire[64:0] T39;
  reg [64:0] R40;
  wire[64:0] T41;
  wire[64:0] mux_data;
  wire[64:0] T42;
  wire[64:0] T43;
  wire[64:0] T44;
  wire[64:0] T45;
  wire[63:0] T46;
  wire[51:0] T47;
  wire[51:0] T48;
  wire[51:0] T49;
  wire[50:0] T50;
  wire[114:0] T51;
  wire[5:0] T52;
  wire[5:0] T121;
  wire[5:0] T122;
  wire[5:0] T123;
  wire[5:0] T124;
  wire[5:0] T125;
  wire[5:0] T126;
  wire[5:0] T127;
  wire[5:0] T128;
  wire[5:0] T129;
  wire[5:0] T130;
  wire[5:0] T131;
  wire[5:0] T132;
  wire[5:0] T133;
  wire[5:0] T134;
  wire[5:0] T135;
  wire[5:0] T136;
  wire[5:0] T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[5:0] T140;
  wire[5:0] T141;
  wire[5:0] T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire[5:0] T146;
  wire[5:0] T147;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[5:0] T150;
  wire[5:0] T151;
  wire[5:0] T152;
  wire[4:0] T153;
  wire[4:0] T154;
  wire[4:0] T155;
  wire[4:0] T156;
  wire[4:0] T157;
  wire[4:0] T158;
  wire[4:0] T159;
  wire[4:0] T160;
  wire[4:0] T161;
  wire[4:0] T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] T166;
  wire[4:0] T167;
  wire[4:0] T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire[3:0] T172;
  wire[3:0] T173;
  wire[3:0] T174;
  wire[3:0] T175;
  wire[3:0] T176;
  wire[2:0] T177;
  wire[2:0] T178;
  wire[2:0] T179;
  wire[2:0] T180;
  wire[1:0] T181;
  wire[1:0] T182;
  wire T183;
  wire[63:0] T54;
  wire[63:0] T55;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T56;
  wire[10:0] T57;
  wire[11:0] T58;
  wire[11:0] T246;
  wire[9:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[1:0] T64;
  wire[11:0] T65;
  wire[11:0] T247;
  wire[10:0] T66;
  wire[10:0] T248;
  wire[1:0] T67;
  wire[11:0] T68;
  wire[11:0] T249;
  wire[11:0] T69;
  wire[11:0] T250;
  wire[11:0] T70;
  wire[11:0] T71;
  wire[11:0] T72;
  wire[2:0] T73;
  wire[2:0] T251;
  wire T74;
  wire T75;
  wire[64:0] T76;
  wire[32:0] T77;
  wire[31:0] T78;
  wire[22:0] T79;
  wire[22:0] T80;
  wire[22:0] T81;
  wire[21:0] T82;
  wire[53:0] T83;
  wire[4:0] T84;
  wire[4:0] T252;
  wire[4:0] T253;
  wire[4:0] T254;
  wire[4:0] T255;
  wire[4:0] T256;
  wire[4:0] T257;
  wire[4:0] T258;
  wire[4:0] T259;
  wire[4:0] T260;
  wire[4:0] T261;
  wire[4:0] T262;
  wire[4:0] T263;
  wire[4:0] T264;
  wire[4:0] T265;
  wire[4:0] T266;
  wire[4:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[3:0] T270;
  wire[3:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[3:0] T274;
  wire[3:0] T275;
  wire[2:0] T276;
  wire[2:0] T277;
  wire[2:0] T278;
  wire[2:0] T279;
  wire[1:0] T280;
  wire[1:0] T281;
  wire T282;
  wire[31:0] T86;
  wire[31:0] T87;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T88;
  wire[7:0] T89;
  wire[8:0] T90;
  wire[8:0] T313;
  wire[6:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[1:0] T96;
  wire[8:0] T97;
  wire[8:0] T314;
  wire[7:0] T98;
  wire[7:0] T315;
  wire[1:0] T99;
  wire[8:0] T100;
  wire[8:0] T316;
  wire[8:0] T101;
  wire[8:0] T317;
  wire[8:0] T102;
  wire[8:0] T103;
  wire[8:0] T104;
  wire[2:0] T105;
  wire[2:0] T318;
  wire T106;
  wire T107;
  wire[64:0] T108;
  reg  R109;
  wire T319;
  wire[32:0] l2s_io_out;
  wire[4:0] l2s_io_exceptionFlags;
  wire[64:0] l2d_io_out;
  wire[4:0] l2d_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R6 = {3{$random}};
    R12 = {1{$random}};
    R21 = {1{$random}};
    R23 = {1{$random}};
    R28 = {1{$random}};
    R32 = {1{$random}};
    R36 = {1{$random}};
    R37 = {1{$random}};
    R38 = {3{$random}};
    R40 = {3{$random}};
    R109 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T110 = R0[1'h1:1'h0];
  assign T1 = io_in_valid ? io_in_bits_rm : R0;
  assign T111 = T2[6'h3f:1'h0];
  assign T2 = longValue;
  assign longValue = T15 ? T14 : T112;
  assign T112 = {T115, T3};
  assign T3 = T11 ? T8 : T113;
  assign T113 = {T114, T4};
  assign T4 = T5;
  assign T5 = R6[5'h1f:1'h0];
  assign T7 = io_in_valid ? io_in_bits_in1 : R6;
  assign T114 = T4[5'h1f];
  assign T8 = T9;
  assign T9 = {1'h0, T10};
  assign T10 = R6[5'h1f:1'h0];
  assign T11 = R12[1'h0];
  assign T13 = io_in_valid ? io_in_bits_typ : R12;
  assign T115 = T116 ? 32'hffffffff : 32'h0;
  assign T116 = T3[6'h20];
  assign T14 = R6;
  assign T15 = R12[1'h1];
  assign T16 = ~ T17;
  assign T17 = R12[1'h0];
  assign T117 = R0[1'h1:1'h0];
  assign T118 = T18[6'h3f:1'h0];
  assign T18 = longValue;
  assign T19 = ~ T20;
  assign T20 = R12[1'h0];
  assign io_out_bits_exc = R21;
  assign T22 = R37 ? R23 : R21;
  assign T24 = R36 ? mux_exc : R23;
  assign mux_exc = T25;
  assign T25 = T34 ? l2d_io_exceptionFlags : T26;
  assign T26 = T27 ? l2s_io_exceptionFlags : 5'h0;
  assign T27 = T30 & R28;
  assign T29 = io_in_valid ? io_in_bits_single : R28;
  assign T30 = 5'h0 == T31;
  assign T31 = R32 & 5'h4;
  assign T33 = io_in_valid ? io_in_bits_cmd : R32;
  assign T34 = T30 & T35;
  assign T35 = R28 ^ 1'h1;
  assign T119 = reset ? 1'h0 : io_in_valid;
  assign T120 = reset ? 1'h0 : R36;
  assign io_out_bits_data = R38;
  assign T39 = R37 ? R40 : R38;
  assign T41 = R36 ? mux_data : R40;
  assign mux_data = T42;
  assign T42 = T34 ? l2d_io_out : T43;
  assign T43 = T27 ? T108 : T44;
  assign T44 = R28 ? T76 : T45;
  assign T45 = {T75, T46};
  assign T46 = {T58, T47};
  assign T47 = T56 ? T49 : T48;
  assign T48 = R6[6'h33:1'h0];
  assign T49 = {T50, 1'h0};
  assign T50 = T51[6'h32:1'h0];
  assign T51 = T48 << T52;
  assign T52 = ~ T121;
  assign T121 = T245 ? 6'h3f : T122;
  assign T122 = T244 ? 6'h3e : T123;
  assign T123 = T243 ? 6'h3d : T124;
  assign T124 = T242 ? 6'h3c : T125;
  assign T125 = T241 ? 6'h3b : T126;
  assign T126 = T240 ? 6'h3a : T127;
  assign T127 = T239 ? 6'h39 : T128;
  assign T128 = T238 ? 6'h38 : T129;
  assign T129 = T237 ? 6'h37 : T130;
  assign T130 = T236 ? 6'h36 : T131;
  assign T131 = T235 ? 6'h35 : T132;
  assign T132 = T234 ? 6'h34 : T133;
  assign T133 = T233 ? 6'h33 : T134;
  assign T134 = T232 ? 6'h32 : T135;
  assign T135 = T231 ? 6'h31 : T136;
  assign T136 = T230 ? 6'h30 : T137;
  assign T137 = T229 ? 6'h2f : T138;
  assign T138 = T228 ? 6'h2e : T139;
  assign T139 = T227 ? 6'h2d : T140;
  assign T140 = T226 ? 6'h2c : T141;
  assign T141 = T225 ? 6'h2b : T142;
  assign T142 = T224 ? 6'h2a : T143;
  assign T143 = T223 ? 6'h29 : T144;
  assign T144 = T222 ? 6'h28 : T145;
  assign T145 = T221 ? 6'h27 : T146;
  assign T146 = T220 ? 6'h26 : T147;
  assign T147 = T219 ? 6'h25 : T148;
  assign T148 = T218 ? 6'h24 : T149;
  assign T149 = T217 ? 6'h23 : T150;
  assign T150 = T216 ? 6'h22 : T151;
  assign T151 = T215 ? 6'h21 : T152;
  assign T152 = T214 ? 6'h20 : T153;
  assign T153 = T213 ? 5'h1f : T154;
  assign T154 = T212 ? 5'h1e : T155;
  assign T155 = T211 ? 5'h1d : T156;
  assign T156 = T210 ? 5'h1c : T157;
  assign T157 = T209 ? 5'h1b : T158;
  assign T158 = T208 ? 5'h1a : T159;
  assign T159 = T207 ? 5'h19 : T160;
  assign T160 = T206 ? 5'h18 : T161;
  assign T161 = T205 ? 5'h17 : T162;
  assign T162 = T204 ? 5'h16 : T163;
  assign T163 = T203 ? 5'h15 : T164;
  assign T164 = T202 ? 5'h14 : T165;
  assign T165 = T201 ? 5'h13 : T166;
  assign T166 = T200 ? 5'h12 : T167;
  assign T167 = T199 ? 5'h11 : T168;
  assign T168 = T198 ? 5'h10 : T169;
  assign T169 = T197 ? 4'hf : T170;
  assign T170 = T196 ? 4'he : T171;
  assign T171 = T195 ? 4'hd : T172;
  assign T172 = T194 ? 4'hc : T173;
  assign T173 = T193 ? 4'hb : T174;
  assign T174 = T192 ? 4'ha : T175;
  assign T175 = T191 ? 4'h9 : T176;
  assign T176 = T190 ? 4'h8 : T177;
  assign T177 = T189 ? 3'h7 : T178;
  assign T178 = T188 ? 3'h6 : T179;
  assign T179 = T187 ? 3'h5 : T180;
  assign T180 = T186 ? 3'h4 : T181;
  assign T181 = T185 ? 2'h3 : T182;
  assign T182 = T184 ? 2'h2 : T183;
  assign T183 = T54[1'h1];
  assign T54 = T55;
  assign T55 = T48 << 4'hc;
  assign T184 = T54[2'h2];
  assign T185 = T54[2'h3];
  assign T186 = T54[3'h4];
  assign T187 = T54[3'h5];
  assign T188 = T54[3'h6];
  assign T189 = T54[3'h7];
  assign T190 = T54[4'h8];
  assign T191 = T54[4'h9];
  assign T192 = T54[4'ha];
  assign T193 = T54[4'hb];
  assign T194 = T54[4'hc];
  assign T195 = T54[4'hd];
  assign T196 = T54[4'he];
  assign T197 = T54[4'hf];
  assign T198 = T54[5'h10];
  assign T199 = T54[5'h11];
  assign T200 = T54[5'h12];
  assign T201 = T54[5'h13];
  assign T202 = T54[5'h14];
  assign T203 = T54[5'h15];
  assign T204 = T54[5'h16];
  assign T205 = T54[5'h17];
  assign T206 = T54[5'h18];
  assign T207 = T54[5'h19];
  assign T208 = T54[5'h1a];
  assign T209 = T54[5'h1b];
  assign T210 = T54[5'h1c];
  assign T211 = T54[5'h1d];
  assign T212 = T54[5'h1e];
  assign T213 = T54[5'h1f];
  assign T214 = T54[6'h20];
  assign T215 = T54[6'h21];
  assign T216 = T54[6'h22];
  assign T217 = T54[6'h23];
  assign T218 = T54[6'h24];
  assign T219 = T54[6'h25];
  assign T220 = T54[6'h26];
  assign T221 = T54[6'h27];
  assign T222 = T54[6'h28];
  assign T223 = T54[6'h29];
  assign T224 = T54[6'h2a];
  assign T225 = T54[6'h2b];
  assign T226 = T54[6'h2c];
  assign T227 = T54[6'h2d];
  assign T228 = T54[6'h2e];
  assign T229 = T54[6'h2f];
  assign T230 = T54[6'h30];
  assign T231 = T54[6'h31];
  assign T232 = T54[6'h32];
  assign T233 = T54[6'h33];
  assign T234 = T54[6'h34];
  assign T235 = T54[6'h35];
  assign T236 = T54[6'h36];
  assign T237 = T54[6'h37];
  assign T238 = T54[6'h38];
  assign T239 = T54[6'h39];
  assign T240 = T54[6'h3a];
  assign T241 = T54[6'h3b];
  assign T242 = T54[6'h3c];
  assign T243 = T54[6'h3d];
  assign T244 = T54[6'h3e];
  assign T245 = T54[6'h3f];
  assign T56 = T57 == 11'h0;
  assign T57 = R6[6'h3e:6'h34];
  assign T58 = T70 | T246;
  assign T246 = {2'h0, T59};
  assign T59 = T60 << 4'h9;
  assign T60 = T63 & T61;
  assign T61 = T62 ^ 1'h1;
  assign T62 = T48 == 52'h0;
  assign T63 = T64 == 2'h3;
  assign T64 = T65[4'hb:4'ha];
  assign T65 = T68 + T247;
  assign T247 = {1'h0, T66};
  assign T66 = 11'h400 | T248;
  assign T248 = {9'h0, T67};
  assign T67 = T56 ? 2'h2 : 2'h1;
  assign T68 = T56 ? T69 : T249;
  assign T249 = {1'h0, T57};
  assign T69 = T250 ^ 12'hfff;
  assign T250 = {6'h0, T52};
  assign T70 = T65 & T71;
  assign T71 = ~ T72;
  assign T72 = T73 << 4'h9;
  assign T73 = 3'h0 - T251;
  assign T251 = {2'h0, T74};
  assign T74 = T56 & T62;
  assign T75 = R6[6'h3f];
  assign T76 = {32'hffffffff, T77};
  assign T77 = {T107, T78};
  assign T78 = {T90, T79};
  assign T79 = T88 ? T81 : T80;
  assign T80 = R6[5'h16:1'h0];
  assign T81 = {T82, 1'h0};
  assign T82 = T83[5'h15:1'h0];
  assign T83 = T80 << T84;
  assign T84 = ~ T252;
  assign T252 = T312 ? 5'h1f : T253;
  assign T253 = T311 ? 5'h1e : T254;
  assign T254 = T310 ? 5'h1d : T255;
  assign T255 = T309 ? 5'h1c : T256;
  assign T256 = T308 ? 5'h1b : T257;
  assign T257 = T307 ? 5'h1a : T258;
  assign T258 = T306 ? 5'h19 : T259;
  assign T259 = T305 ? 5'h18 : T260;
  assign T260 = T304 ? 5'h17 : T261;
  assign T261 = T303 ? 5'h16 : T262;
  assign T262 = T302 ? 5'h15 : T263;
  assign T263 = T301 ? 5'h14 : T264;
  assign T264 = T300 ? 5'h13 : T265;
  assign T265 = T299 ? 5'h12 : T266;
  assign T266 = T298 ? 5'h11 : T267;
  assign T267 = T297 ? 5'h10 : T268;
  assign T268 = T296 ? 4'hf : T269;
  assign T269 = T295 ? 4'he : T270;
  assign T270 = T294 ? 4'hd : T271;
  assign T271 = T293 ? 4'hc : T272;
  assign T272 = T292 ? 4'hb : T273;
  assign T273 = T291 ? 4'ha : T274;
  assign T274 = T290 ? 4'h9 : T275;
  assign T275 = T289 ? 4'h8 : T276;
  assign T276 = T288 ? 3'h7 : T277;
  assign T277 = T287 ? 3'h6 : T278;
  assign T278 = T286 ? 3'h5 : T279;
  assign T279 = T285 ? 3'h4 : T280;
  assign T280 = T284 ? 2'h3 : T281;
  assign T281 = T283 ? 2'h2 : T282;
  assign T282 = T86[1'h1];
  assign T86 = T87;
  assign T87 = T80 << 4'h9;
  assign T283 = T86[2'h2];
  assign T284 = T86[2'h3];
  assign T285 = T86[3'h4];
  assign T286 = T86[3'h5];
  assign T287 = T86[3'h6];
  assign T288 = T86[3'h7];
  assign T289 = T86[4'h8];
  assign T290 = T86[4'h9];
  assign T291 = T86[4'ha];
  assign T292 = T86[4'hb];
  assign T293 = T86[4'hc];
  assign T294 = T86[4'hd];
  assign T295 = T86[4'he];
  assign T296 = T86[4'hf];
  assign T297 = T86[5'h10];
  assign T298 = T86[5'h11];
  assign T299 = T86[5'h12];
  assign T300 = T86[5'h13];
  assign T301 = T86[5'h14];
  assign T302 = T86[5'h15];
  assign T303 = T86[5'h16];
  assign T304 = T86[5'h17];
  assign T305 = T86[5'h18];
  assign T306 = T86[5'h19];
  assign T307 = T86[5'h1a];
  assign T308 = T86[5'h1b];
  assign T309 = T86[5'h1c];
  assign T310 = T86[5'h1d];
  assign T311 = T86[5'h1e];
  assign T312 = T86[5'h1f];
  assign T88 = T89 == 8'h0;
  assign T89 = R6[5'h1e:5'h17];
  assign T90 = T102 | T313;
  assign T313 = {2'h0, T91};
  assign T91 = T92 << 3'h6;
  assign T92 = T95 & T93;
  assign T93 = T94 ^ 1'h1;
  assign T94 = T80 == 23'h0;
  assign T95 = T96 == 2'h3;
  assign T96 = T97[4'h8:3'h7];
  assign T97 = T100 + T314;
  assign T314 = {1'h0, T98};
  assign T98 = 8'h80 | T315;
  assign T315 = {6'h0, T99};
  assign T99 = T88 ? 2'h2 : 2'h1;
  assign T100 = T88 ? T101 : T316;
  assign T316 = {1'h0, T89};
  assign T101 = T317 ^ 9'h1ff;
  assign T317 = {4'h0, T84};
  assign T102 = T97 & T103;
  assign T103 = ~ T104;
  assign T104 = T105 << 3'h6;
  assign T105 = 3'h0 - T318;
  assign T318 = {2'h0, T106};
  assign T106 = T88 & T94;
  assign T107 = R6[5'h1f];
  assign T108 = {32'hffffffff, l2s_io_out};
  assign io_out_valid = R109;
  assign T319 = reset ? 1'h0 : R37;
  INToRecFN_0 l2s(
       .io_signedIn( T19 ),
       .io_in( T118 ),
       .io_roundingMode( T117 ),
       .io_out( l2s_io_out ),
       .io_exceptionFlags( l2s_io_exceptionFlags )
  );
  INToRecFN_1 l2d(
       .io_signedIn( T16 ),
       .io_in( T111 ),
       .io_roundingMode( T110 ),
       .io_out( l2d_io_out ),
       .io_exceptionFlags( l2d_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      R0 <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      R6 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R12 <= io_in_bits_typ;
    end
    if(R37) begin
      R21 <= R23;
    end
    if(R36) begin
      R23 <= mux_exc;
    end
    if(io_in_valid) begin
      R28 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R32 <= io_in_bits_cmd;
    end
    if(reset) begin
      R36 <= 1'h0;
    end else begin
      R36 <= io_in_valid;
    end
    if(reset) begin
      R37 <= 1'h0;
    end else begin
      R37 <= R36;
    end
    if(R37) begin
      R38 <= R40;
    end
    if(R36) begin
      R40 <= mux_data;
    end
    if(reset) begin
      R109 <= 1'h0;
    end else begin
      R109 <= R37;
    end
  end
endmodule

module RoundRawFNToRecFN(
    input  io_invalidExc,
    input  io_infiniteExc,
    input  io_in_sign,
    input  io_in_isNaN,
    input  io_in_isInf,
    input  io_in_isZero,
    input [9:0] io_in_sExp,
    input [26:0] io_in_sig,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire anyRound;
  wire anyRoundExtra;
  wire[26:0] T4;
  wire[26:0] T127;
  wire[25:0] T5;
  wire[26:0] roundMask;
  wire[24:0] T6;
  wire[24:0] T128;
  wire doShiftSigDown1;
  wire[24:0] T7;
  wire[24:0] T8;
  wire[8:0] T9;
  wire T10;
  wire[8:0] T11;
  wire[24:0] T12;
  wire[512:0] T13;
  wire[8:0] T14;
  wire[8:0] T15;
  wire[7:0] T16;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[6:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[5:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[7:0] T26;
  wire[3:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T129;
  wire[3:0] T30;
  wire[7:0] T31;
  wire[7:0] T130;
  wire[5:0] T32;
  wire[7:0] T33;
  wire[7:0] T131;
  wire[6:0] T34;
  wire[15:0] T35;
  wire[15:0] T36;
  wire[15:0] T37;
  wire[14:0] T38;
  wire[15:0] T39;
  wire[15:0] T40;
  wire[15:0] T41;
  wire[13:0] T42;
  wire[15:0] T43;
  wire[15:0] T44;
  wire[15:0] T45;
  wire[11:0] T46;
  wire[15:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[7:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire[15:0] T132;
  wire[7:0] T53;
  wire[15:0] T54;
  wire[15:0] T133;
  wire[11:0] T55;
  wire[15:0] T56;
  wire[15:0] T134;
  wire[13:0] T57;
  wire[15:0] T58;
  wire[15:0] T135;
  wire[14:0] T59;
  wire[24:0] T60;
  wire[24:0] T136;
  wire T61;
  wire roundPosBit;
  wire[26:0] T62;
  wire[26:0] roundPosMask;
  wire[26:0] T137;
  wire[25:0] T63;
  wire[25:0] T64;
  wire commonCase;
  wire T65;
  wire T66;
  wire T67;
  wire notNaN_isSpecialInfOut;
  wire T68;
  wire isNaNOut;
  wire underflow;
  wire common_underflow;
  wire T69;
  wire[8:0] T70;
  wire overflow;
  wire common_overflow;
  wire[2:0] T71;
  wire[9:0] sRoundedExp;
  wire[9:0] T138;
  wire[2:0] T72;
  wire[2:0] T73;
  wire[1:0] T74;
  wire[25:0] roundedSig;
  wire[25:0] T139;
  wire[24:0] T75;
  wire[26:0] T76;
  wire[26:0] T77;
  wire[25:0] T78;
  wire[25:0] T79;
  wire[25:0] T80;
  wire[25:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire roundingMode_nearest_even;
  wire[25:0] T140;
  wire[24:0] T85;
  wire[24:0] T86;
  wire[26:0] T87;
  wire T88;
  wire T89;
  wire roundMagUp;
  wire T90;
  wire T91;
  wire roundingMode_max;
  wire T92;
  wire roundingMode_min;
  wire T93;
  wire[6:0] T141;
  wire T142;
  wire[1:0] T94;
  wire[32:0] T95;
  wire[31:0] T96;
  wire[22:0] fractOut;
  wire[22:0] T97;
  wire[22:0] T143;
  wire pegMaxFiniteMagOut;
  wire T98;
  wire overflow_roundMagUp;
  wire T99;
  wire[22:0] T100;
  wire[22:0] common_fractOut;
  wire[22:0] T101;
  wire[22:0] T102;
  wire[22:0] T103;
  wire T104;
  wire common_totalUnderflow;
  wire[8:0] expOut;
  wire[8:0] T105;
  wire[8:0] T106;
  wire[8:0] T107;
  wire notNaN_isInfOut;
  wire T108;
  wire[8:0] T109;
  wire[8:0] T110;
  wire[8:0] T111;
  wire[8:0] T112;
  wire pegMinNonzeroMagOut;
  wire T113;
  wire[8:0] T114;
  wire[8:0] T115;
  wire[8:0] T116;
  wire[8:0] T117;
  wire[8:0] T118;
  wire[8:0] T119;
  wire[8:0] T120;
  wire[8:0] T121;
  wire[8:0] T122;
  wire[8:0] T123;
  wire[8:0] T124;
  wire[8:0] T125;
  wire T126;
  wire[8:0] common_expOut;
  wire signOut;


  assign io_exceptionFlags = T0;
  assign T0 = {T94, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 27'h0;
  assign T4 = io_in_sig & T127;
  assign T127 = {1'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = {T6, 2'h3};
  assign T6 = T7 | T128;
  assign T128 = {24'h0, doShiftSigDown1};
  assign doShiftSigDown1 = io_in_sig[5'h1a];
  assign T7 = T60 | T8;
  assign T8 = {T35, T9};
  assign T9 = {T16, T10};
  assign T10 = T11[4'h8];
  assign T11 = T12[5'h18:5'h10];
  assign T12 = T13[8'h82:7'h6a];
  assign T13 = $signed(513'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T14;
  assign T14 = ~ T15;
  assign T15 = io_in_sExp[4'h8:1'h0];
  assign T16 = T33 | T17;
  assign T17 = T18 & 8'haa;
  assign T18 = T19 << 1'h1;
  assign T19 = T20[3'h6:1'h0];
  assign T20 = T31 | T21;
  assign T21 = T22 & 8'hcc;
  assign T22 = T23 << 2'h2;
  assign T23 = T24[3'h5:1'h0];
  assign T24 = T29 | T25;
  assign T25 = T26 & 8'hf0;
  assign T26 = T27 << 3'h4;
  assign T27 = T28[2'h3:1'h0];
  assign T28 = T11[3'h7:1'h0];
  assign T29 = T129 & 8'hf;
  assign T129 = {4'h0, T30};
  assign T30 = T28 >> 3'h4;
  assign T31 = T130 & 8'h33;
  assign T130 = {2'h0, T32};
  assign T32 = T24 >> 2'h2;
  assign T33 = T131 & 8'h55;
  assign T131 = {1'h0, T34};
  assign T34 = T20 >> 1'h1;
  assign T35 = T58 | T36;
  assign T36 = T37 & 16'haaaa;
  assign T37 = T38 << 1'h1;
  assign T38 = T39[4'he:1'h0];
  assign T39 = T56 | T40;
  assign T40 = T41 & 16'hcccc;
  assign T41 = T42 << 2'h2;
  assign T42 = T43[4'hd:1'h0];
  assign T43 = T54 | T44;
  assign T44 = T45 & 16'hf0f0;
  assign T45 = T46 << 3'h4;
  assign T46 = T47[4'hb:1'h0];
  assign T47 = T52 | T48;
  assign T48 = T49 & 16'hff00;
  assign T49 = T50 << 4'h8;
  assign T50 = T51[3'h7:1'h0];
  assign T51 = T12[4'hf:1'h0];
  assign T52 = T132 & 16'hff;
  assign T132 = {8'h0, T53};
  assign T53 = T51 >> 4'h8;
  assign T54 = T133 & 16'hf0f;
  assign T133 = {4'h0, T55};
  assign T55 = T47 >> 3'h4;
  assign T56 = T134 & 16'h3333;
  assign T134 = {2'h0, T57};
  assign T57 = T43 >> 2'h2;
  assign T58 = T135 & 16'h5555;
  assign T135 = {1'h0, T59};
  assign T59 = T39 >> 1'h1;
  assign T60 = 25'h0 - T136;
  assign T136 = {24'h0, T61};
  assign T61 = $signed(io_in_sExp) < $signed(1'h0);
  assign roundPosBit = T62 != 27'h0;
  assign T62 = io_in_sig & roundPosMask;
  assign roundPosMask = T137 & roundMask;
  assign T137 = {1'h0, T63};
  assign T63 = ~ T64;
  assign T64 = roundMask >> 1'h1;
  assign commonCase = T66 & T65;
  assign T65 = io_in_isZero ^ 1'h1;
  assign T66 = T68 & T67;
  assign T67 = notNaN_isSpecialInfOut ^ 1'h1;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T68 = isNaNOut ^ 1'h1;
  assign isNaNOut = io_invalidExc | io_in_isNaN;
  assign underflow = commonCase & common_underflow;
  assign common_underflow = anyRound & T69;
  assign T69 = $signed(io_in_sExp) < $signed(T70);
  assign T70 = doShiftSigDown1 ? 9'h81 : 9'h82;
  assign overflow = commonCase & common_overflow;
  assign common_overflow = $signed(3'h3) <= $signed(T71);
  assign T71 = $signed(sRoundedExp) >>> 3'h7;
  assign sRoundedExp = io_in_sExp + T138;
  assign T138 = {T141, T72};
  assign T72 = T73;
  assign T73 = {1'h0, T74};
  assign T74 = roundedSig >> 5'h18;
  assign roundedSig = T88 ? T78 : T139;
  assign T139 = {1'h0, T75};
  assign T75 = T76 >> 2'h2;
  assign T76 = io_in_sig & T77;
  assign T77 = ~ roundMask;
  assign T78 = T140 & T79;
  assign T79 = ~ T80;
  assign T80 = T82 ? T81 : 26'h0;
  assign T81 = roundMask >> 1'h1;
  assign T82 = T84 & T83;
  assign T83 = anyRoundExtra ^ 1'h1;
  assign T84 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T140 = {1'h0, T85};
  assign T85 = T86 + 25'h1;
  assign T86 = T87 >> 2'h2;
  assign T87 = io_in_sig | roundMask;
  assign T88 = T93 | T89;
  assign T89 = roundMagUp & anyRound;
  assign roundMagUp = T92 | T90;
  assign T90 = roundingMode_max & T91;
  assign T91 = io_in_sign ^ 1'h1;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign T92 = roundingMode_min & io_in_sign;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign T93 = roundingMode_nearest_even & roundPosBit;
  assign T141 = T142 ? 7'h7f : 7'h0;
  assign T142 = T72[2'h2];
  assign T94 = {io_invalidExc, io_infiniteExc};
  assign io_out = T95;
  assign T95 = {signOut, T96};
  assign T96 = {expOut, fractOut};
  assign fractOut = T100 | T97;
  assign T97 = 23'h0 - T143;
  assign T143 = {22'h0, pegMaxFiniteMagOut};
  assign pegMaxFiniteMagOut = T99 & T98;
  assign T98 = overflow_roundMagUp ^ 1'h1;
  assign overflow_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign T99 = commonCase & overflow;
  assign T100 = T104 ? T103 : common_fractOut;
  assign common_fractOut = doShiftSigDown1 ? T102 : T101;
  assign T101 = roundedSig[5'h16:1'h0];
  assign T102 = roundedSig[5'h17:1'h1];
  assign T103 = isNaNOut ? 23'h400000 : 23'h0;
  assign T104 = common_totalUnderflow | isNaNOut;
  assign common_totalUnderflow = $signed(sRoundedExp) < $signed(8'h6b);
  assign expOut = T106 | T105;
  assign T105 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T106 = T109 | T107;
  assign T107 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T108;
  assign T108 = overflow & overflow_roundMagUp;
  assign T109 = T111 | T110;
  assign T110 = pegMaxFiniteMagOut ? 9'h17f : 9'h0;
  assign T111 = T114 | T112;
  assign T112 = pegMinNonzeroMagOut ? 9'h6b : 9'h0;
  assign pegMinNonzeroMagOut = T113 & roundMagUp;
  assign T113 = commonCase & common_totalUnderflow;
  assign T114 = T117 & T115;
  assign T115 = ~ T116;
  assign T116 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T117 = T120 & T118;
  assign T118 = ~ T119;
  assign T119 = pegMaxFiniteMagOut ? 9'h80 : 9'h0;
  assign T120 = T123 & T121;
  assign T121 = ~ T122;
  assign T122 = pegMinNonzeroMagOut ? 9'h194 : 9'h0;
  assign T123 = common_expOut & T124;
  assign T124 = ~ T125;
  assign T125 = T126 ? 9'h1c0 : 9'h0;
  assign T126 = io_in_isZero | common_totalUnderflow;
  assign common_expOut = sRoundedExp[4'h8:1'h0];
  assign signOut = isNaNOut ? 1'h0 : io_in_sign;
endmodule

module RecFNToRecFN_1(
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[26:0] outRawFloat_sig;
  wire[26:0] T0;
  wire T1;
  wire[29:0] T2;
  wire[55:0] T3;
  wire[55:0] T4;
  wire[53:0] T5;
  wire[51:0] T6;
  wire[25:0] T7;
  wire[9:0] outRawFloat_sExp;
  wire[9:0] T8;
  wire[9:0] T9;
  wire[8:0] T10;
  wire[8:0] T11;
  wire[12:0] T12;
  wire[12:0] T13;
  wire[12:0] T14;
  wire[12:0] T15;
  wire[11:0] T16;
  wire T17;
  wire[2:0] T18;
  wire T19;
  wire outRawFloat_isZero;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire outRawFloat_isInf;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire outRawFloat_isNaN;
  wire T29;
  wire T30;
  wire T31;
  wire outRawFloat_sign;
  wire T32;
  wire T33;
  wire invalidExc;
  wire T34;
  wire T35;
  wire[32:0] RoundRawFNToRecFN_io_out;
  wire[4:0] RoundRawFNToRecFN_io_exceptionFlags;


  assign outRawFloat_sig = T0;
  assign T0 = {T7, T1};
  assign T1 = T2 != 30'h0;
  assign T2 = T3[5'h1d:1'h0];
  assign T3 = T4;
  assign T4 = {2'h1, T5};
  assign T5 = {T6, 2'h0};
  assign T6 = io_in[6'h33:1'h0];
  assign T7 = T3[6'h37:5'h1e];
  assign outRawFloat_sExp = T8;
  assign T8 = T9;
  assign T9 = {T19, T10};
  assign T10 = T17 ? 9'h1fc : T11;
  assign T11 = T12[4'h8:1'h0];
  assign T12 = T13 + 13'h1900;
  assign T13 = T14;
  assign T14 = T15;
  assign T15 = {1'h0, T16};
  assign T16 = io_in[6'h3f:6'h34];
  assign T17 = T18 != 3'h0;
  assign T18 = T12[4'hb:4'h9];
  assign T19 = $signed(T12) < $signed(1'h0);
  assign outRawFloat_isZero = T20;
  assign T20 = T21;
  assign T21 = T22 == 3'h0;
  assign T22 = T16[4'hb:4'h9];
  assign outRawFloat_isInf = T23;
  assign T23 = T24;
  assign T24 = T27 & T25;
  assign T25 = T26 ^ 1'h1;
  assign T26 = T16[4'h9];
  assign T27 = T28 == 2'h3;
  assign T28 = T16[4'hb:4'ha];
  assign outRawFloat_isNaN = T29;
  assign T29 = T30;
  assign T30 = T27 & T31;
  assign T31 = T16[4'h9];
  assign outRawFloat_sign = T32;
  assign T32 = T33;
  assign T33 = io_in[7'h40];
  assign invalidExc = outRawFloat_isNaN & T34;
  assign T34 = T35 ^ 1'h1;
  assign T35 = outRawFloat_sig[5'h18];
  assign io_exceptionFlags = RoundRawFNToRecFN_io_exceptionFlags;
  assign io_out = RoundRawFNToRecFN_io_out;
  RoundRawFNToRecFN RoundRawFNToRecFN(
       .io_invalidExc( invalidExc ),
       .io_infiniteExc( 1'h0 ),
       .io_in_sign( outRawFloat_sign ),
       .io_in_isNaN( outRawFloat_isNaN ),
       .io_in_isInf( outRawFloat_isInf ),
       .io_in_isZero( outRawFloat_isZero ),
       .io_in_sExp( outRawFloat_sExp ),
       .io_in_sig( outRawFloat_sig ),
       .io_roundingMode( io_roundingMode ),
       .io_out( RoundRawFNToRecFN_io_out ),
       .io_exceptionFlags( RoundRawFNToRecFN_io_exceptionFlags )
  );
endmodule

module FPToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap12,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_div,
    input  io_in_bits_sqrt,
    input  io_in_bits_round,
    input  io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc,
    input  io_lt
);

  wire[1:0] T73;
  reg [2:0] R0;
  wire[2:0] T1;
  reg [64:0] R2;
  wire[64:0] T3;
  wire[1:0] T74;
  wire[32:0] T75;
  reg [4:0] R4;
  wire[4:0] T5;
  wire[4:0] mux_exc;
  wire[4:0] T6;
  wire[4:0] T7;
  wire[4:0] T8;
  wire[4:0] minmax_exc;
  wire T9;
  wire issnan2;
  wire T10;
  wire T11;
  wire T12;
  reg [64:0] R13;
  wire[64:0] T14;
  wire T15;
  reg  R16;
  wire T17;
  wire isnan2;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire issnan1;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire isnan1;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire[2:0] T29;
  wire isSgnj;
  wire[4:0] T30;
  reg [4:0] R31;
  wire[4:0] T32;
  wire T33;
  wire T34;
  wire[4:0] T35;
  wire T36;
  wire T37;
  reg  R38;
  wire T76;
  reg [64:0] R39;
  wire[64:0] T40;
  wire[64:0] mux_data;
  wire[64:0] T41;
  wire[64:0] T42;
  wire[64:0] T43;
  wire[64:0] fsgnj;
  wire[32:0] T44;
  wire[31:0] T45;
  wire sign_s;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[31:0] T55;
  wire[30:0] T56;
  wire sign_d;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire isLHS;
  wire T68;
  wire T69;
  wire T70;
  wire isMax;
  wire[64:0] T71;
  reg  R72;
  wire T77;
  wire[64:0] s2d_io_out;
  wire[4:0] s2d_io_exceptionFlags;
  wire[32:0] d2s_io_out;
  wire[4:0] d2s_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R2 = {3{$random}};
    R4 = {1{$random}};
    R13 = {3{$random}};
    R16 = {1{$random}};
    R31 = {1{$random}};
    R38 = {1{$random}};
    R39 = {3{$random}};
    R72 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T73 = R0[1'h1:1'h0];
  assign T1 = io_in_valid ? io_in_bits_rm : R0;
  assign T3 = io_in_valid ? io_in_bits_in1 : R2;
  assign T74 = R0[1'h1:1'h0];
  assign T75 = R2[6'h20:1'h0];
  assign io_out_bits_exc = R4;
  assign T5 = R38 ? mux_exc : R4;
  assign mux_exc = T6;
  assign T6 = T36 ? s2d_io_exceptionFlags : T7;
  assign T7 = T33 ? d2s_io_exceptionFlags : T8;
  assign T8 = isSgnj ? 5'h0 : minmax_exc;
  assign minmax_exc = {T9, 4'h0};
  assign T9 = issnan1 | issnan2;
  assign issnan2 = isnan2 & T10;
  assign T10 = ~ T11;
  assign T11 = R16 ? T15 : T12;
  assign T12 = R13[6'h33];
  assign T14 = io_in_valid ? io_in_bits_in2 : R13;
  assign T15 = R13[5'h16];
  assign T17 = io_in_valid ? io_in_bits_single : R16;
  assign isnan2 = R16 ? T20 : T18;
  assign T18 = T19 == 3'h7;
  assign T19 = R13[6'h3f:6'h3d];
  assign T20 = T21 == 3'h7;
  assign T21 = R13[5'h1f:5'h1d];
  assign issnan1 = isnan1 & T22;
  assign T22 = ~ T23;
  assign T23 = R16 ? T25 : T24;
  assign T24 = R2[6'h33];
  assign T25 = R2[5'h16];
  assign isnan1 = R16 ? T28 : T26;
  assign T26 = T27 == 3'h7;
  assign T27 = R2[6'h3f:6'h3d];
  assign T28 = T29 == 3'h7;
  assign T29 = R2[5'h1f:5'h1d];
  assign isSgnj = 5'h4 == T30;
  assign T30 = R31 & 5'h5;
  assign T32 = io_in_valid ? io_in_bits_cmd : R31;
  assign T33 = T34 & R16;
  assign T34 = 5'h0 == T35;
  assign T35 = R31 & 5'h4;
  assign T36 = T34 & T37;
  assign T37 = R16 ^ 1'h1;
  assign T76 = reset ? 1'h0 : io_in_valid;
  assign io_out_bits_data = R39;
  assign T40 = R38 ? mux_data : R39;
  assign mux_data = T41;
  assign T41 = T36 ? s2d_io_out : T42;
  assign T42 = T33 ? T71 : T43;
  assign T43 = T67 ? fsgnj : R13;
  assign fsgnj = {T55, T44};
  assign T44 = {sign_s, T45};
  assign T45 = R2[5'h1f:1'h0];
  assign sign_s = T49 ^ T46;
  assign T46 = T48 & T47;
  assign T47 = R13[6'h20];
  assign T48 = R16 & isSgnj;
  assign T49 = T52 ? T51 : T50;
  assign T50 = R0[1'h0];
  assign T51 = R2[6'h20];
  assign T52 = T54 | T53;
  assign T53 = T48 ^ 1'h1;
  assign T54 = R0[1'h1];
  assign T55 = {sign_d, T56};
  assign T56 = R2[6'h3f:6'h21];
  assign sign_d = T61 ^ T57;
  assign T57 = T59 & T58;
  assign T58 = R13[7'h40];
  assign T59 = T60 & isSgnj;
  assign T60 = R16 ^ 1'h1;
  assign T61 = T64 ? T63 : T62;
  assign T62 = R0[1'h0];
  assign T63 = R2[7'h40];
  assign T64 = T66 | T65;
  assign T65 = T59 ^ 1'h1;
  assign T66 = R0[1'h1];
  assign T67 = isSgnj | isLHS;
  assign isLHS = isnan2 | T68;
  assign T68 = T70 & T69;
  assign T69 = isnan1 ^ 1'h1;
  assign T70 = isMax != io_lt;
  assign isMax = R0[1'h0];
  assign T71 = {32'hffffffff, d2s_io_out};
  assign io_out_valid = R72;
  assign T77 = reset ? 1'h0 : R38;
  RecFNToRecFN s2d(
       .io_in( T75 ),
       .io_roundingMode( T74 ),
       .io_out( s2d_io_out ),
       .io_exceptionFlags( s2d_io_exceptionFlags )
  );
  RecFNToRecFN_1 d2s(
       .io_in( R2 ),
       .io_roundingMode( T73 ),
       .io_out( d2s_io_out ),
       .io_exceptionFlags( d2s_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      R0 <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      R2 <= io_in_bits_in1;
    end
    if(R38) begin
      R4 <= mux_exc;
    end
    if(io_in_valid) begin
      R13 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      R16 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R31 <= io_in_bits_cmd;
    end
    if(reset) begin
      R38 <= 1'h0;
    end else begin
      R38 <= io_in_valid;
    end
    if(R38) begin
      R39 <= mux_data;
    end
    if(reset) begin
      R72 <= 1'h0;
    end else begin
      R72 <= R38;
    end
  end
endmodule

module DivSqrtRecF64_mulAddZ31(input clk, input reset,
    output io_inReady_div,
    output io_inReady_sqrt,
    input  io_inValid,
    input  io_sqrtOp,
    input [64:0] io_a,
    input [64:0] io_b,
    input [1:0] io_roundingMode,
    output io_outValid_div,
    output io_outValid_sqrt,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags,
    output[3:0] io_usingMulAdd,
    output io_latchMulAddA_0,
    output[53:0] io_mulAddA_0,
    output io_latchMulAddB_0,
    output[53:0] io_mulAddB_0,
    output[104:0] io_mulAddC_2,
    input [104:0] io_mulAddResult_3
);

  wire[104:0] T0;
  wire[104:0] T885;
  wire[55:0] T1;
  wire[55:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  reg  extraT_E;
  wire T6;
  wire T7;
  wire[53:0] sigT_C1;
  wire[53:0] zComplSigT_C1;
  wire[53:0] T8;
  wire[53:0] T9;
  wire[53:0] T10;
  wire[52:0] T11;
  wire[52:0] T12;
  wire T13;
  wire E_C1_div;
  wire T14;
  wire cyc_C1_div;
  wire T15;
  reg  sqrtOp_PC;
  wire T16;
  wire T17;
  reg  sqrtOp_PB;
  wire T18;
  wire T19;
  reg  sqrtOp_PA;
  wire T20;
  wire entering_PA;
  wire T21;
  wire T22;
  wire T23;
  wire ready_PB;
  wire T24;
  wire valid_leaving_PB;
  wire ready_PC;
  wire T25;
  wire valid_leaving_PC;
  wire cyc_E1;
  wire T26;
  reg [2:0] cycleNum_E;
  wire[2:0] T886;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire normalCase_PC;
  wire T33;
  wire T34;
  wire isZeroB_PC;
  reg [2:0] specialCodeB_PC;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] specialCodeB_S;
  wire[11:0] expB_S;
  reg [2:0] specialCodeB_PB;
  wire[2:0] T37;
  wire[2:0] T38;
  reg [2:0] specialCodeB_PA;
  wire[2:0] T39;
  wire T40;
  wire T41;
  wire isZeroA_PC;
  reg [2:0] specialCodeA_PC;
  wire[2:0] T42;
  wire[2:0] T43;
  wire[2:0] specialCodeA_S;
  wire[11:0] expA_S;
  reg [2:0] specialCodeA_PB;
  wire[2:0] T44;
  wire[2:0] T45;
  reg [2:0] specialCodeA_PA;
  wire[2:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire isSpecialB_PC;
  wire[1:0] T51;
  wire T52;
  wire isSpecialA_PC;
  wire[1:0] T53;
  wire T54;
  wire T55;
  reg  sign_PC;
  wire T56;
  wire T57;
  wire sign_S;
  wire T58;
  wire signA_S;
  wire signB_S;
  reg  sign_PB;
  wire T59;
  wire T60;
  reg  sign_PA;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  reg  valid_PC;
  wire T887;
  wire T66;
  wire T67;
  wire leaving_PC;
  wire T68;
  wire cyc_C3;
  wire T69;
  reg [2:0] cycleNum_C;
  wire[2:0] T888;
  wire[2:0] T70;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire cyc_B1;
  wire T74;
  reg [3:0] cycleNum_B;
  wire[3:0] T889;
  wire[3:0] T75;
  wire[3:0] T76;
  wire[3:0] T77;
  wire[3:0] T78;
  wire cyc_A1;
  reg [2:0] cycleNum_A;
  wire[2:0] T890;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire T83;
  wire[2:0] T84;
  wire[2:0] T85;
  wire cyc_A7_sqrt;
  wire normalCase_S_sqrt;
  wire T86;
  wire T87;
  wire T88;
  wire isZeroB_S;
  wire T89;
  wire isSpecialB_S;
  wire[1:0] T90;
  wire cyc_S_sqrt;
  wire T91;
  wire[2:0] T891;
  wire[1:0] T92;
  wire cyc_A4_div;
  wire normalCase_S_div;
  wire T93;
  wire T94;
  wire T95;
  wire isZeroA_S;
  wire T96;
  wire T97;
  wire T98;
  wire isSpecialA_S;
  wire[1:0] T99;
  wire cyc_S_div;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire normalCase_PB;
  wire T108;
  wire T109;
  wire isZeroB_PB;
  wire T110;
  wire T111;
  wire isZeroA_PB;
  wire T112;
  wire T113;
  wire isSpecialB_PB;
  wire[1:0] T114;
  wire T115;
  wire isSpecialA_PB;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire cyc_S;
  wire entering_PA_normalCase;
  reg  valid_PA;
  wire T892;
  wire T123;
  wire T124;
  wire leaving_PA;
  wire T125;
  wire valid_leaving_PA;
  wire valid_normalCase_leaving_PA;
  wire cyc_B7_sqrt;
  wire T126;
  wire cyc_B4_div;
  wire T127;
  wire T128;
  wire T129;
  wire cyc_B4;
  wire T130;
  wire normalCase_PA;
  wire T131;
  wire T132;
  wire isZeroB_PA;
  wire T133;
  wire T134;
  wire isZeroA_PA;
  wire T135;
  wire T136;
  wire isSpecialB_PA;
  wire[1:0] T137;
  wire T138;
  wire isSpecialA_PA;
  wire[1:0] T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire entering_PB;
  wire entering_PB_S;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire leaving_PB;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire normalCase_S;
  reg  valid_PB;
  wire T893;
  wire T154;
  wire T155;
  wire entering_PC;
  wire entering_PC_S;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[53:0] T162;
  wire[53:0] T163;
  wire[53:0] T164;
  wire T165;
  wire cyc_C1_sqrt;
  wire T166;
  wire T167;
  wire cyc_C1;
  wire T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire T171;
  wire[52:0] sigB_PC;
  wire[51:0] T172;
  reg [50:0] fractB_other_PC;
  wire[50:0] T173;
  reg [50:0] fractB_other_PB;
  wire[50:0] T174;
  reg [50:0] fractB_other_PA;
  wire[50:0] T175;
  wire[50:0] T176;
  wire[51:0] fractB_S;
  wire entering_PB_normalCase;
  wire T177;
  wire entering_PC_normalCase;
  wire T178;
  reg  fractB_51_PC;
  wire T179;
  wire T180;
  wire T181;
  reg  fractB_51_PB;
  wire T182;
  wire T183;
  wire T184;
  reg  fractB_51_PA;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  reg [13:0] exp_PC;
  wire[13:0] T193;
  reg [13:0] exp_PB;
  wire[13:0] T194;
  reg [13:0] exp_PA;
  wire[13:0] T195;
  wire[13:0] T196;
  wire[13:0] T197;
  wire[13:0] T198;
  wire[10:0] T199;
  wire[10:0] T200;
  wire[2:0] T201;
  wire[2:0] T894;
  wire T202;
  wire[13:0] T895;
  wire[13:0] T896;
  wire cyc_E3_sqrt;
  wire cyc_E3;
  wire T203;
  wire[104:0] T204;
  wire[104:0] T897;
  wire[53:0] T205;
  wire[53:0] T206;
  reg  fractA_0_PC;
  wire T207;
  reg  fractA_0_PB;
  wire T208;
  wire T209;
  reg [50:0] fractA_other_PA;
  wire[50:0] T210;
  wire[50:0] T211;
  wire[51:0] fractA_S;
  wire T212;
  wire T213;
  reg  E_E_div;
  wire T214;
  wire cyc_E3_div;
  wire T215;
  wire[104:0] T216;
  wire[104:0] T217;
  wire[104:0] T218;
  reg [57:0] sigXN_C;
  wire[57:0] T219;
  wire[57:0] sigXNU_B3_CX;
  wire[57:0] T220;
  wire T221;
  wire cyc_C3_sqrt;
  wire T222;
  wire cyc_C5_div;
  wire T223;
  wire cyc_C5;
  wire T224;
  wire cyc_C6_sqrt;
  wire T225;
  wire cyc_C2;
  wire T226;
  wire cyc_C4_sqrt;
  wire cyc_C4;
  wire T227;
  wire[104:0] T228;
  wire[104:0] T898;
  wire[103:0] T229;
  wire[103:0] T230;
  reg [57:0] sigX1_B;
  wire[57:0] T231;
  wire cyc_B3;
  wire T232;
  wire[104:0] T233;
  wire[104:0] T234;
  wire[53:0] T235;
  wire[53:0] T899;
  wire[52:0] T236;
  wire[52:0] T900;
  wire[32:0] T237;
  reg [32:0] sqrSigma1_C;
  wire[32:0] T238;
  wire[32:0] sqrSigma1_B1;
  wire[52:0] T239;
  wire[52:0] T901;
  wire[29:0] T240;
  wire[29:0] T241;
  wire[52:0] T242;
  wire[52:0] T902;
  wire[45:0] zSigma1_B4;
  wire[45:0] T243;
  wire[45:0] T244;
  wire[45:0] T245;
  wire[52:0] T246;
  wire[52:0] T247;
  wire[52:0] T248;
  reg [16:0] ER1_B_sqrt;
  wire[16:0] T249;
  wire[16:0] ER1_A1_sqrt;
  wire[16:0] T903;
  wire[15:0] r1_A1;
  wire[14:0] fractR1_A1;
  wire[15:0] T250;
  wire[15:0] T251;
  wire[24:0] mulAdd9Out_A;
  wire[17:0] T252;
  wire[18:0] loMulAdd9Out_A;
  wire[18:0] T253;
  wire[17:0] T254;
  wire[24:0] mulAdd9C_A;
  wire[24:0] T904;
  wire[23:0] T255;
  wire[23:0] T256;
  reg [8:0] fractR0_A;
  wire[8:0] T257;
  wire[8:0] T258;
  wire[8:0] zFractR0_A4_div;
  wire[13:0] T259;
  wire[13:0] T260;
  wire[24:0] T261;
  wire T262;
  wire T263;
  wire[8:0] zFractR0_A6_sqrt;
  wire[14:0] T264;
  wire[14:0] T265;
  wire[24:0] T266;
  wire T267;
  wire T268;
  wire cyc_A6_sqrt;
  wire T269;
  wire cyc_A1_div;
  wire T270;
  wire[24:0] T271;
  wire[24:0] T272;
  wire[24:0] T273;
  wire[24:0] T905;
  wire[20:0] T274;
  wire[20:0] T275;
  reg [20:0] partNegSigma0_A;
  wire[20:0] T276;
  wire[20:0] T277;
  wire[24:0] T278;
  wire[24:0] T906;
  wire[15:0] T279;
  wire cyc_A4_sqrt;
  wire T280;
  wire cyc_A3;
  wire T281;
  wire cyc_A2;
  wire cyc_A3_sqrt;
  wire[20:0] T282;
  wire[20:0] T283;
  wire[20:0] T284;
  wire[20:0] T285;
  wire[52:0] sigB_PA;
  wire[51:0] T286;
  wire T287;
  wire cyc_A3_div;
  wire T288;
  wire T289;
  wire T290;
  reg [9:0] hiSqrR0_A_sqrt;
  wire[9:0] T907;
  wire[15:0] T291;
  wire[15:0] T908;
  wire[15:0] T292;
  wire[25:0] sqrR0_A5_sqrt;
  wire[25:0] T909;
  wire[25:0] T293;
  wire T294;
  wire cyc_A5_sqrt;
  wire[20:0] T295;
  wire[20:0] T910;
  wire[10:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire[20:0] T300;
  wire[20:0] T911;
  wire[19:0] T301;
  wire[19:0] T302;
  wire[19:0] T912;
  wire[18:0] T303;
  wire[20:0] T304;
  wire[20:0] T305;
  wire[19:0] T306;
  wire[7:0] T307;
  wire[7:0] T913;
  wire[11:0] zComplFractK0_A4_div;
  wire[11:0] T308;
  wire zLinPiece_7_A4_div;
  wire T309;
  wire[2:0] T310;
  wire[11:0] T311;
  wire[11:0] T312;
  wire zLinPiece_6_A4_div;
  wire T313;
  wire[2:0] T314;
  wire[11:0] T315;
  wire[11:0] T316;
  wire zLinPiece_5_A4_div;
  wire T317;
  wire[2:0] T318;
  wire[11:0] T319;
  wire[11:0] T320;
  wire zLinPiece_4_A4_div;
  wire T321;
  wire[2:0] T322;
  wire[11:0] T323;
  wire[11:0] T324;
  wire zLinPiece_3_A4_div;
  wire T325;
  wire[2:0] T326;
  wire[11:0] T327;
  wire[11:0] T328;
  wire zLinPiece_2_A4_div;
  wire T329;
  wire[2:0] T330;
  wire[11:0] T331;
  wire[11:0] T332;
  wire zLinPiece_1_A4_div;
  wire T333;
  wire[2:0] T334;
  wire[11:0] T335;
  wire zLinPiece_0_A4_div;
  wire T336;
  wire[2:0] T337;
  wire[20:0] T914;
  wire[19:0] T338;
  wire[19:0] T339;
  wire[18:0] T340;
  wire[5:0] T341;
  wire[5:0] T915;
  wire[12:0] zComplFractK0_A6_sqrt;
  wire[12:0] T342;
  wire zQuadPiece_3_A6_sqrt;
  wire T343;
  wire T344;
  wire T345;
  wire[12:0] T346;
  wire[12:0] T347;
  wire zQuadPiece_2_A6_sqrt;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire[12:0] T352;
  wire[12:0] T353;
  wire zQuadPiece_1_A6_sqrt;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire[12:0] T358;
  wire zQuadPiece_0_A6_sqrt;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire[19:0] T364;
  wire[9:0] T365;
  wire[9:0] T916;
  wire[9:0] zComplK1_A7_sqrt;
  wire[9:0] T366;
  wire zQuadPiece_3_A7_sqrt;
  wire T367;
  wire T368;
  wire T369;
  wire[9:0] T370;
  wire[9:0] T371;
  wire zQuadPiece_2_A7_sqrt;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[9:0] T376;
  wire[9:0] T377;
  wire zQuadPiece_1_A7_sqrt;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[9:0] T382;
  wire zQuadPiece_0_A7_sqrt;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[18:0] T917;
  wire[17:0] T388;
  wire[8:0] mulAdd9B_A;
  wire[8:0] T389;
  reg [8:0] nextMulAdd9B_A;
  wire[8:0] T390;
  wire[8:0] T391;
  wire[8:0] T392;
  wire[8:0] T393;
  wire[7:0] T394;
  wire[8:0] T395;
  wire[8:0] T396;
  wire[8:0] T397;
  wire[8:0] T398;
  wire[8:0] T399;
  wire[8:0] T400;
  wire[8:0] T401;
  wire[8:0] T402;
  wire[8:0] T403;
  wire[51:0] zFractB_A7_sqrt;
  wire T404;
  wire T405;
  wire cyc_A4;
  wire T406;
  wire T407;
  wire T408;
  wire[8:0] T409;
  wire[8:0] T410;
  wire[8:0] zK1_A4_div;
  wire[8:0] T411;
  wire[8:0] T412;
  wire[8:0] T413;
  wire[8:0] T414;
  wire[8:0] T415;
  wire[8:0] T416;
  wire[8:0] T417;
  wire[8:0] T418;
  wire[8:0] T419;
  wire[8:0] T420;
  wire[8:0] T421;
  wire[8:0] T422;
  wire[8:0] T423;
  wire[8:0] T424;
  wire[8:0] mulAdd9A_A;
  wire[8:0] T425;
  reg [8:0] nextMulAdd9A_A;
  wire[8:0] T918;
  wire[13:0] T426;
  wire[13:0] T919;
  wire[13:0] T427;
  wire[13:0] T920;
  wire[8:0] zSigma0_A2;
  wire[22:0] T428;
  wire[22:0] T429;
  wire[24:0] T430;
  wire T431;
  wire T432;
  wire[13:0] T433;
  wire[13:0] T921;
  wire[8:0] T434;
  wire[8:0] T435;
  wire T436;
  wire[13:0] T437;
  wire[13:0] T922;
  wire[8:0] T438;
  wire[51:0] zFractB_A4_div;
  wire[13:0] T439;
  wire[13:0] T923;
  wire[8:0] T440;
  wire[8:0] T441;
  wire[13:0] T442;
  wire[13:0] T924;
  wire[13:0] T443;
  wire[13:0] T444;
  wire[24:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[8:0] T452;
  wire[8:0] zK2_A7_sqrt;
  wire[8:0] T453;
  wire[8:0] T454;
  wire[8:0] T455;
  wire[8:0] T456;
  wire[8:0] T457;
  wire[8:0] T458;
  wire[8:0] T459;
  wire[6:0] T460;
  wire[6:0] T461;
  wire[6:0] T462;
  wire[6:0] T463;
  wire T464;
  wire[15:0] T925;
  wire[14:0] T465;
  wire[16:0] T466;
  wire T467;
  wire cyc_A1_sqrt;
  wire cyc_B6_sqrt;
  wire T468;
  wire T469;
  wire cyc_B6;
  wire T470;
  wire[52:0] T926;
  wire[51:0] T471;
  wire[51:0] T927;
  wire[50:0] T472;
  wire[50:0] T473;
  reg [31:0] ESqrR1_B_sqrt;
  wire[31:0] T474;
  wire[31:0] ESqrR1_B8_sqrt;
  wire cyc_B8_sqrt;
  wire T475;
  wire[51:0] T476;
  wire[51:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[53:0] T484;
  wire[53:0] zComplSigT_C1_sqrt;
  wire[53:0] T485;
  wire[53:0] T486;
  wire[53:0] T487;
  wire[53:0] T928;
  wire[52:0] T488;
  wire[52:0] T489;
  wire[52:0] T490;
  wire[52:0] T929;
  wire[45:0] T491;
  wire[45:0] T492;
  reg [30:0] u_C_sqrt;
  wire[30:0] T493;
  wire[30:0] T494;
  wire cyc_C5_sqrt;
  wire[52:0] T495;
  wire[52:0] T930;
  wire[45:0] T496;
  wire[45:0] T497;
  wire[32:0] T498;
  wire cyc_C4_div;
  wire T499;
  wire[52:0] T500;
  wire[52:0] T931;
  wire[45:0] T501;
  wire[45:0] T502;
  wire T503;
  wire[52:0] T504;
  wire[52:0] T932;
  wire[33:0] T505;
  wire[52:0] T506;
  wire[52:0] T507;
  wire[52:0] sigA_PA;
  wire[51:0] T508;
  reg  fractA_51_PA;
  wire T509;
  wire T510;
  wire cyc_B6_div;
  wire T511;
  wire T512;
  wire T513;
  wire[52:0] T514;
  wire[52:0] T515;
  wire T516;
  wire[52:0] T517;
  wire[52:0] T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[3:0] T526;
  wire[1:0] T527;
  wire T528;
  wire cyc_B2_sqrt;
  wire T529;
  wire cyc_B2;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire cyc_B1_sqrt;
  wire T535;
  wire T536;
  wire cyc_B3_sqrt;
  wire T537;
  wire T538;
  wire T539;
  wire cyc_B5;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire T545;
  wire T546;
  wire T547;
  wire cyc_B1_div;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire cyc_B4_sqrt;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire cyc_B9_sqrt;
  wire T558;
  wire T559;
  wire cyc_A2_div;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire cyc_B2_div;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire cyc_B5_sqrt;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire cyc_B10_sqrt;
  wire T574;
  wire T575;
  wire T576;
  wire[4:0] T577;
  wire[2:0] T578;
  wire[1:0] T579;
  wire inexact_E1;
  wire T580;
  wire inexactY_E1;
  wire anyRoundExtra_E1;
  wire T581;
  wire all1sHiRoundExtraT_E;
  wire[52:0] T582;
  wire[52:0] T933;
  wire[51:0] T583;
  wire[52:0] roundMask_E;
  wire[20:0] T584;
  wire[4:0] T585;
  wire T586;
  wire[4:0] T587;
  wire[20:0] T588;
  wire[52:0] T589;
  wire[8192:0] T590;
  wire[12:0] T591;
  wire[12:0] posExpX_E;
  wire[13:0] sExpX_E;
  wire[13:0] T934;
  wire[12:0] T592;
  wire[12:0] T593;
  wire[12:0] T594;
  wire[13:0] T595;
  wire[13:0] T596;
  wire[13:0] expP1_PC;
  wire[13:0] T597;
  wire[12:0] T598;
  wire[13:0] T599;
  wire[12:0] T600;
  wire[13:0] expP2_PC;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire[13:0] T605;
  wire T606;
  wire T607;
  wire[3:0] T608;
  wire[1:0] T609;
  wire T610;
  wire[1:0] T611;
  wire[3:0] T612;
  wire T613;
  wire[1:0] T614;
  wire T615;
  wire[1:0] T616;
  wire T617;
  wire[15:0] T618;
  wire[15:0] T619;
  wire[15:0] T620;
  wire[14:0] T621;
  wire[15:0] T622;
  wire[15:0] T623;
  wire[15:0] T624;
  wire[13:0] T625;
  wire[15:0] T626;
  wire[15:0] T627;
  wire[15:0] T628;
  wire[11:0] T629;
  wire[15:0] T630;
  wire[15:0] T631;
  wire[15:0] T632;
  wire[7:0] T633;
  wire[15:0] T634;
  wire[15:0] T635;
  wire[15:0] T935;
  wire[7:0] T636;
  wire[15:0] T637;
  wire[15:0] T936;
  wire[11:0] T638;
  wire[15:0] T639;
  wire[15:0] T937;
  wire[13:0] T640;
  wire[15:0] T641;
  wire[15:0] T938;
  wire[14:0] T642;
  wire[31:0] T643;
  wire[31:0] T644;
  wire[31:0] T645;
  wire[30:0] T646;
  wire[31:0] T647;
  wire[31:0] T648;
  wire[31:0] T649;
  wire[29:0] T650;
  wire[31:0] T651;
  wire[31:0] T652;
  wire[31:0] T653;
  wire[27:0] T654;
  wire[31:0] T655;
  wire[31:0] T656;
  wire[31:0] T657;
  wire[23:0] T658;
  wire[31:0] T659;
  wire[31:0] T660;
  wire[31:0] T661;
  wire[15:0] T662;
  wire[31:0] T663;
  wire[31:0] T664;
  wire[31:0] T939;
  wire[15:0] T665;
  wire[31:0] T666;
  wire[31:0] T940;
  wire[23:0] T667;
  wire[31:0] T668;
  wire[31:0] T941;
  wire[27:0] T669;
  wire[31:0] T670;
  wire[31:0] T942;
  wire[29:0] T671;
  wire[31:0] T672;
  wire[31:0] T943;
  wire[30:0] T673;
  wire[52:0] T674;
  reg [52:0] sigT_E;
  wire[52:0] T675;
  wire[52:0] T676;
  wire T677;
  wire T678;
  wire T679;
  reg  isZeroRemT_E;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[55:0] remT_E2;
  wire T685;
  wire T686;
  wire[53:0] T687;
  wire cyc_E2;
  wire T688;
  wire hiRoundPosBit_E1;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire trueLtX_E1;
  reg  isNegRemT_E;
  wire T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire hiRoundPosBitT_E;
  wire[52:0] T701;
  wire[52:0] T702;
  wire[53:0] incrPosMask_E;
  wire[53:0] T703;
  wire[53:0] T704;
  wire[53:0] T705;
  wire T706;
  wire underflow_E1;
  wire underflowY_E1;
  wire T707;
  wire T708;
  wire totalUnderflowY_E1;
  wire T709;
  wire[12:0] T710;
  wire[13:0] sExpY_E1;
  wire[13:0] T944;
  wire[12:0] T711;
  wire[12:0] T712;
  wire[12:0] T713;
  wire T714;
  wire T715;
  wire[53:0] sigY_E1;
  wire[53:0] T716;
  wire[53:0] roundEvenMask_E1;
  wire T717;
  wire T718;
  wire T719;
  wire roundingMode_near_even_PC;
  reg [1:0] roundingMode_PC;
  wire[1:0] T720;
  wire[1:0] T721;
  reg [1:0] roundingMode_PB;
  wire[1:0] T722;
  wire[1:0] T723;
  reg [1:0] roundingMode_PA;
  wire[1:0] T724;
  wire[53:0] T725;
  wire[53:0] sigY0_E;
  wire[53:0] T726;
  wire[52:0] T727;
  wire[53:0] sigAdjT_E;
  wire[53:0] T945;
  wire roundMagUp_PC;
  wire roundingMode_max_PC;
  wire roundingMode_min_PC;
  wire[53:0] T728;
  wire[53:0] T946;
  wire[53:0] sigY1_E;
  wire[53:0] T729;
  wire[53:0] T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire all1sHiRoundT_E;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire roundMagDown_PC;
  wire T758;
  wire T759;
  wire[13:0] T760;
  wire[13:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[13:0] T767;
  wire[13:0] T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire[13:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire overflow_E1;
  wire overflowY_E1;
  wire T777;
  wire[2:0] T778;
  wire T779;
  wire T780;
  wire[1:0] T781;
  wire infinity_PC;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire invalid_PC;
  wire notSigNaN_invalid_PC;
  wire T787;
  wire T788;
  wire isInfB_PC;
  wire T789;
  wire T790;
  wire isInfA_PC;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire isNaNB_PC;
  wire T798;
  wire T799;
  wire isSigNaNB_PC;
  wire T800;
  wire T801;
  wire isSigNaNA_PC;
  wire T802;
  reg  fractA_51_PC;
  wire T803;
  wire T804;
  wire T805;
  reg  fractA_51_PB;
  wire T806;
  wire T807;
  wire T808;
  wire isNaNA_PC;
  wire T809;
  wire T810;
  wire[64:0] T811;
  wire[63:0] T812;
  wire[51:0] fractOut_E1;
  wire[51:0] T813;
  wire[51:0] T947;
  wire pegMaxFiniteMagOut_E1;
  wire T814;
  wire overflowY_roundMagUp_PC;
  wire[51:0] T815;
  wire[51:0] fractY_E1;
  wire[51:0] T816;
  wire isNaNOut_PC;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire notSpecial_isZeroOut_E1;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire[11:0] expOut_E1;
  wire[11:0] T826;
  wire[11:0] T827;
  wire[11:0] T828;
  wire notNaN_isInfOut_E1;
  wire T829;
  wire T830;
  wire T831;
  wire[11:0] T832;
  wire[11:0] T833;
  wire[11:0] T834;
  wire[11:0] T835;
  wire pegMinFiniteMagOut_E1;
  wire T836;
  wire[11:0] T837;
  wire[11:0] T838;
  wire[11:0] T839;
  wire[11:0] T840;
  wire[11:0] T841;
  wire[11:0] T842;
  wire[11:0] T843;
  wire[11:0] T844;
  wire[11:0] T845;
  wire[11:0] T846;
  wire[11:0] T847;
  wire[11:0] T848;
  wire[11:0] expY_E1;
  wire signOut_PC;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire ready_PA;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    extraT_E = {1{$random}};
    sqrtOp_PC = {1{$random}};
    sqrtOp_PB = {1{$random}};
    sqrtOp_PA = {1{$random}};
    cycleNum_E = {1{$random}};
    specialCodeB_PC = {1{$random}};
    specialCodeB_PB = {1{$random}};
    specialCodeB_PA = {1{$random}};
    specialCodeA_PC = {1{$random}};
    specialCodeA_PB = {1{$random}};
    specialCodeA_PA = {1{$random}};
    sign_PC = {1{$random}};
    sign_PB = {1{$random}};
    sign_PA = {1{$random}};
    valid_PC = {1{$random}};
    cycleNum_C = {1{$random}};
    cycleNum_B = {1{$random}};
    cycleNum_A = {1{$random}};
    valid_PA = {1{$random}};
    valid_PB = {1{$random}};
    fractB_other_PC = {2{$random}};
    fractB_other_PB = {2{$random}};
    fractB_other_PA = {2{$random}};
    fractB_51_PC = {1{$random}};
    fractB_51_PB = {1{$random}};
    fractB_51_PA = {1{$random}};
    exp_PC = {1{$random}};
    exp_PB = {1{$random}};
    exp_PA = {1{$random}};
    fractA_0_PC = {1{$random}};
    fractA_0_PB = {1{$random}};
    fractA_other_PA = {2{$random}};
    E_E_div = {1{$random}};
    sigXN_C = {2{$random}};
    sigX1_B = {2{$random}};
    sqrSigma1_C = {2{$random}};
    ER1_B_sqrt = {1{$random}};
    fractR0_A = {1{$random}};
    partNegSigma0_A = {1{$random}};
    hiSqrR0_A_sqrt = {1{$random}};
    nextMulAdd9B_A = {1{$random}};
    nextMulAdd9A_A = {1{$random}};
    ESqrR1_B_sqrt = {1{$random}};
    u_C_sqrt = {1{$random}};
    fractA_51_PA = {1{$random}};
    sigT_E = {2{$random}};
    isZeroRemT_E = {1{$random}};
    isNegRemT_E = {1{$random}};
    roundingMode_PC = {1{$random}};
    roundingMode_PB = {1{$random}};
    roundingMode_PA = {1{$random}};
    fractA_51_PC = {1{$random}};
    fractA_51_PB = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_mulAddC_2 = T0;
  assign T0 = T204 | T885;
  assign T885 = {49'h0, T1};
  assign T1 = cyc_E3_sqrt ? T2 : 56'h0;
  assign T2 = T3 << 6'h36;
  assign T3 = T169 ^ T4;
  assign T4 = {T5, 1'h0};
  assign T5 = extraT_E ^ 1'h1;
  assign T6 = cyc_C1 ? T7 : extraT_E;
  assign T7 = sigT_C1[1'h0];
  assign sigT_C1 = ~ zComplSigT_C1;
  assign zComplSigT_C1 = T8;
  assign T8 = T162 | T9;
  assign T9 = T13 ? T10 : 54'h0;
  assign T10 = {1'h0, T11};
  assign T11 = ~ T12;
  assign T12 = io_mulAddResult_3[7'h66:6'h32];
  assign T13 = cyc_C1_div & E_C1_div;
  assign E_C1_div = T14 ^ 1'h1;
  assign T14 = io_mulAddResult_3[7'h68];
  assign cyc_C1_div = cyc_C1 & T15;
  assign T15 = sqrtOp_PC ^ 1'h1;
  assign T16 = entering_PC ? T17 : sqrtOp_PC;
  assign T17 = valid_PB ? sqrtOp_PB : io_sqrtOp;
  assign T18 = entering_PB ? T19 : sqrtOp_PB;
  assign T19 = valid_PA ? sqrtOp_PA : io_sqrtOp;
  assign T20 = entering_PA ? io_sqrtOp : sqrtOp_PA;
  assign entering_PA = entering_PA_normalCase | T21;
  assign T21 = cyc_S & T22;
  assign T22 = valid_PA | T23;
  assign T23 = ready_PB ^ 1'h1;
  assign ready_PB = T24;
  assign T24 = T122 | valid_leaving_PB;
  assign valid_leaving_PB = normalCase_PB ? cyc_C3 : ready_PC;
  assign ready_PC = T25;
  assign T25 = T65 | valid_leaving_PC;
  assign valid_leaving_PC = T32 | cyc_E1;
  assign cyc_E1 = T26;
  assign T26 = cycleNum_E == 3'h1;
  assign T886 = reset ? 3'h0 : T27;
  assign T27 = T30 ? T28 : cycleNum_E;
  assign T28 = cyc_C1 ? 3'h4 : T29;
  assign T29 = cycleNum_E - 3'h1;
  assign T30 = cyc_C1 | T31;
  assign T31 = cycleNum_E != 3'h0;
  assign T32 = normalCase_PC ^ 1'h1;
  assign normalCase_PC = sqrtOp_PC ? T54 : T33;
  assign T33 = T40 & T34;
  assign T34 = isZeroB_PC ^ 1'h1;
  assign isZeroB_PC = specialCodeB_PC == 3'h0;
  assign T35 = entering_PC ? T36 : specialCodeB_PC;
  assign T36 = valid_PB ? specialCodeB_PB : specialCodeB_S;
  assign specialCodeB_S = expB_S[4'hb:4'h9];
  assign expB_S = io_b[6'h3f:6'h34];
  assign T37 = entering_PB ? T38 : specialCodeB_PB;
  assign T38 = valid_PA ? specialCodeB_PA : specialCodeB_S;
  assign T39 = entering_PA ? specialCodeB_S : specialCodeB_PA;
  assign T40 = T49 & T41;
  assign T41 = isZeroA_PC ^ 1'h1;
  assign isZeroA_PC = specialCodeA_PC == 3'h0;
  assign T42 = entering_PC ? T43 : specialCodeA_PC;
  assign T43 = valid_PB ? specialCodeA_PB : specialCodeA_S;
  assign specialCodeA_S = expA_S[4'hb:4'h9];
  assign expA_S = io_a[6'h3f:6'h34];
  assign T44 = entering_PB ? T45 : specialCodeA_PB;
  assign T45 = valid_PA ? specialCodeA_PA : specialCodeA_S;
  assign T46 = T47 ? specialCodeA_S : specialCodeA_PA;
  assign T47 = entering_PA & T48;
  assign T48 = io_sqrtOp ^ 1'h1;
  assign T49 = T52 & T50;
  assign T50 = isSpecialB_PC ^ 1'h1;
  assign isSpecialB_PC = T51 == 2'h3;
  assign T51 = specialCodeB_PC[2'h2:1'h1];
  assign T52 = isSpecialA_PC ^ 1'h1;
  assign isSpecialA_PC = T53 == 2'h3;
  assign T53 = specialCodeA_PC[2'h2:1'h1];
  assign T54 = T62 & T55;
  assign T55 = sign_PC ^ 1'h1;
  assign T56 = entering_PC ? T57 : sign_PC;
  assign T57 = valid_PB ? sign_PB : sign_S;
  assign sign_S = io_sqrtOp ? signB_S : T58;
  assign T58 = signA_S ^ signB_S;
  assign signA_S = io_a[7'h40];
  assign signB_S = io_b[7'h40];
  assign T59 = entering_PB ? T60 : sign_PB;
  assign T60 = valid_PA ? sign_PA : sign_S;
  assign T61 = entering_PA ? sign_S : sign_PA;
  assign T62 = T64 & T63;
  assign T63 = isZeroB_PC ^ 1'h1;
  assign T64 = isSpecialB_PC ^ 1'h1;
  assign T65 = valid_PC ^ 1'h1;
  assign T887 = reset ? 1'h0 : T66;
  assign T66 = T67 ? entering_PC : valid_PC;
  assign T67 = entering_PC | leaving_PC;
  assign leaving_PC = T68;
  assign T68 = valid_PC & valid_leaving_PC;
  assign cyc_C3 = T69;
  assign T69 = cycleNum_C == 3'h3;
  assign T888 = reset ? 3'h0 : T70;
  assign T70 = T106 ? T71 : cycleNum_C;
  assign T71 = cyc_B1 ? T73 : T72;
  assign T72 = cycleNum_C - 3'h1;
  assign T73 = sqrtOp_PB ? 3'h6 : 3'h5;
  assign cyc_B1 = T74;
  assign T74 = cycleNum_B == 4'h1;
  assign T889 = reset ? 4'h0 : T75;
  assign T75 = T104 ? T76 : cycleNum_B;
  assign T76 = cyc_A1 ? T78 : T77;
  assign T77 = cycleNum_B - 4'h1;
  assign T78 = sqrtOp_PA ? 4'ha : 4'h6;
  assign cyc_A1 = cycleNum_A == 3'h1;
  assign T890 = reset ? 3'h0 : T79;
  assign T79 = T102 ? T80 : cycleNum_A;
  assign T80 = T84 | T81;
  assign T81 = T83 ? T82 : 3'h0;
  assign T82 = cycleNum_A - 3'h1;
  assign T83 = entering_PA_normalCase ^ 1'h1;
  assign T84 = T891 | T85;
  assign T85 = cyc_A7_sqrt ? 3'h6 : 3'h0;
  assign cyc_A7_sqrt = cyc_S_sqrt & normalCase_S_sqrt;
  assign normalCase_S_sqrt = T87 & T86;
  assign T86 = signB_S ^ 1'h1;
  assign T87 = T89 & T88;
  assign T88 = isZeroB_S ^ 1'h1;
  assign isZeroB_S = specialCodeB_S == 3'h0;
  assign T89 = isSpecialB_S ^ 1'h1;
  assign isSpecialB_S = T90 == 2'h3;
  assign T90 = specialCodeB_S[2'h2:1'h1];
  assign cyc_S_sqrt = T91 & io_sqrtOp;
  assign T91 = io_inReady_sqrt & io_inValid;
  assign T891 = {1'h0, T92};
  assign T92 = cyc_A4_div ? 2'h3 : 2'h0;
  assign cyc_A4_div = cyc_S_div & normalCase_S_div;
  assign normalCase_S_div = T94 & T93;
  assign T93 = isZeroB_S ^ 1'h1;
  assign T94 = T96 & T95;
  assign T95 = isZeroA_S ^ 1'h1;
  assign isZeroA_S = specialCodeA_S == 3'h0;
  assign T96 = T98 & T97;
  assign T97 = isSpecialB_S ^ 1'h1;
  assign T98 = isSpecialA_S ^ 1'h1;
  assign isSpecialA_S = T99 == 2'h3;
  assign T99 = specialCodeA_S[2'h2:1'h1];
  assign cyc_S_div = T101 & T100;
  assign T100 = io_sqrtOp ^ 1'h1;
  assign T101 = io_inReady_div & io_inValid;
  assign T102 = entering_PA_normalCase | T103;
  assign T103 = cycleNum_A != 3'h0;
  assign T104 = cyc_A1 | T105;
  assign T105 = cycleNum_B != 4'h0;
  assign T106 = cyc_B1 | T107;
  assign T107 = cycleNum_C != 3'h0;
  assign normalCase_PB = sqrtOp_PB ? T117 : T108;
  assign T108 = T110 & T109;
  assign T109 = isZeroB_PB ^ 1'h1;
  assign isZeroB_PB = specialCodeB_PB == 3'h0;
  assign T110 = T112 & T111;
  assign T111 = isZeroA_PB ^ 1'h1;
  assign isZeroA_PB = specialCodeA_PB == 3'h0;
  assign T112 = T115 & T113;
  assign T113 = isSpecialB_PB ^ 1'h1;
  assign isSpecialB_PB = T114 == 2'h3;
  assign T114 = specialCodeB_PB[2'h2:1'h1];
  assign T115 = isSpecialA_PB ^ 1'h1;
  assign isSpecialA_PB = T116 == 2'h3;
  assign T116 = specialCodeA_PB[2'h2:1'h1];
  assign T117 = T119 & T118;
  assign T118 = sign_PB ^ 1'h1;
  assign T119 = T121 & T120;
  assign T120 = isZeroB_PB ^ 1'h1;
  assign T121 = isSpecialB_PB ^ 1'h1;
  assign T122 = valid_PB ^ 1'h1;
  assign cyc_S = cyc_S_div | cyc_S_sqrt;
  assign entering_PA_normalCase = cyc_A4_div | cyc_A7_sqrt;
  assign T892 = reset ? 1'h0 : T123;
  assign T123 = T124 ? entering_PA : valid_PA;
  assign T124 = entering_PA | leaving_PA;
  assign leaving_PA = T125;
  assign T125 = valid_PA & valid_leaving_PA;
  assign valid_leaving_PA = normalCase_PA ? valid_normalCase_leaving_PA : ready_PB;
  assign valid_normalCase_leaving_PA = cyc_B4_div | cyc_B7_sqrt;
  assign cyc_B7_sqrt = T126;
  assign T126 = cycleNum_B == 4'h7;
  assign cyc_B4_div = T127;
  assign T127 = T129 & T128;
  assign T128 = sqrtOp_PA ^ 1'h1;
  assign T129 = cyc_B4 & valid_PA;
  assign cyc_B4 = T130;
  assign T130 = cycleNum_B == 4'h4;
  assign normalCase_PA = sqrtOp_PA ? T140 : T131;
  assign T131 = T133 & T132;
  assign T132 = isZeroB_PA ^ 1'h1;
  assign isZeroB_PA = specialCodeB_PA == 3'h0;
  assign T133 = T135 & T134;
  assign T134 = isZeroA_PA ^ 1'h1;
  assign isZeroA_PA = specialCodeA_PA == 3'h0;
  assign T135 = T138 & T136;
  assign T136 = isSpecialB_PA ^ 1'h1;
  assign isSpecialB_PA = T137 == 2'h3;
  assign T137 = specialCodeB_PA[2'h2:1'h1];
  assign T138 = isSpecialA_PA ^ 1'h1;
  assign isSpecialA_PA = T139 == 2'h3;
  assign T139 = specialCodeA_PA[2'h2:1'h1];
  assign T140 = T142 & T141;
  assign T141 = sign_PA ^ 1'h1;
  assign T142 = T144 & T143;
  assign T143 = isZeroB_PA ^ 1'h1;
  assign T144 = isSpecialB_PA ^ 1'h1;
  assign entering_PB = entering_PB_S | leaving_PA;
  assign entering_PB_S = T150 & T145;
  assign T145 = leaving_PB | T146;
  assign T146 = T148 & T147;
  assign T147 = ready_PC ^ 1'h1;
  assign T148 = valid_PB ^ 1'h1;
  assign leaving_PB = T149;
  assign T149 = valid_PB & valid_leaving_PB;
  assign T150 = T152 & T151;
  assign T151 = valid_PA ^ 1'h1;
  assign T152 = cyc_S & T153;
  assign T153 = normalCase_S ^ 1'h1;
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div;
  assign T893 = reset ? 1'h0 : T154;
  assign T154 = T155 ? entering_PB : valid_PB;
  assign T155 = entering_PB | leaving_PB;
  assign entering_PC = entering_PC_S | leaving_PB;
  assign entering_PC_S = T156 & ready_PC;
  assign T156 = T158 & T157;
  assign T157 = valid_PB ^ 1'h1;
  assign T158 = T160 & T159;
  assign T159 = valid_PA ^ 1'h1;
  assign T160 = cyc_S & T161;
  assign T161 = normalCase_S ^ 1'h1;
  assign T162 = T165 ? T163 : 54'h0;
  assign T163 = ~ T164;
  assign T164 = io_mulAddResult_3[7'h68:6'h33];
  assign T165 = T166 | cyc_C1_sqrt;
  assign cyc_C1_sqrt = cyc_C1 & sqrtOp_PC;
  assign T166 = cyc_C1_div & T167;
  assign T167 = E_C1_div ^ 1'h1;
  assign cyc_C1 = T168;
  assign T168 = cycleNum_C == 3'h1;
  assign T169 = T192 ? T190 : T170;
  assign T170 = {T187, T171};
  assign T171 = sigB_PC[1'h0];
  assign sigB_PC = {1'h1, T172};
  assign T172 = {fractB_51_PC, fractB_other_PC};
  assign T173 = entering_PC_normalCase ? fractB_other_PB : fractB_other_PC;
  assign T174 = entering_PB_normalCase ? fractB_other_PA : fractB_other_PB;
  assign T175 = entering_PA_normalCase ? T176 : fractB_other_PA;
  assign T176 = fractB_S[6'h32:1'h0];
  assign fractB_S = io_b[6'h33:1'h0];
  assign entering_PB_normalCase = T177 & valid_normalCase_leaving_PA;
  assign T177 = valid_PA & normalCase_PA;
  assign entering_PC_normalCase = T178 & cyc_C3;
  assign T178 = valid_PB & normalCase_PB;
  assign T179 = entering_PC ? T180 : fractB_51_PC;
  assign T180 = valid_PB ? fractB_51_PB : T181;
  assign T181 = fractB_S[6'h33];
  assign T182 = entering_PB ? T183 : fractB_51_PB;
  assign T183 = valid_PA ? fractB_51_PA : T184;
  assign T184 = fractB_S[6'h33];
  assign T185 = entering_PA ? T186 : fractB_51_PA;
  assign T186 = fractB_S[6'h33];
  assign T187 = T189 ^ T188;
  assign T188 = sigB_PC[1'h0];
  assign T189 = sigB_PC[1'h1];
  assign T190 = {T191, 1'h0};
  assign T191 = sigB_PC[1'h0];
  assign T192 = exp_PC[1'h0];
  assign T193 = entering_PC_normalCase ? exp_PB : exp_PC;
  assign T194 = entering_PB_normalCase ? exp_PA : exp_PB;
  assign T195 = entering_PA_normalCase ? T196 : exp_PA;
  assign T196 = io_sqrtOp ? T896 : T197;
  assign T197 = T895 + T198;
  assign T198 = {T201, T199};
  assign T199 = ~ T200;
  assign T200 = expB_S[4'ha:1'h0];
  assign T201 = 3'h0 - T894;
  assign T894 = {2'h0, T202};
  assign T202 = expB_S[4'hb];
  assign T895 = {2'h0, expA_S};
  assign T896 = {2'h0, expB_S};
  assign cyc_E3_sqrt = cyc_E3 & sqrtOp_PC;
  assign cyc_E3 = T203;
  assign T203 = cycleNum_E == 3'h3;
  assign T204 = T216 | T897;
  assign T897 = {51'h0, T205};
  assign T205 = T212 ? T206 : 54'h0;
  assign T206 = fractA_0_PC << 6'h35;
  assign T207 = entering_PC_normalCase ? fractA_0_PB : fractA_0_PC;
  assign T208 = entering_PB_normalCase ? T209 : fractA_0_PB;
  assign T209 = fractA_other_PA[1'h0];
  assign T210 = cyc_A4_div ? T211 : fractA_other_PA;
  assign T211 = fractA_S[6'h32:1'h0];
  assign fractA_S = io_a[6'h33:1'h0];
  assign T212 = cyc_E3_div & T213;
  assign T213 = E_E_div ^ 1'h1;
  assign T214 = cyc_C1 ? E_C1_div : E_E_div;
  assign cyc_E3_div = cyc_E3 & T215;
  assign T215 = sqrtOp_PC ^ 1'h1;
  assign T216 = T228 | T217;
  assign T217 = T225 ? T218 : 105'h0;
  assign T218 = sigXN_C << 6'h2f;
  assign T219 = T221 ? sigXNU_B3_CX : sigXN_C;
  assign sigXNU_B3_CX = T220;
  assign T220 = io_mulAddResult_3[7'h68:6'h2f];
  assign T221 = T222 | cyc_C3_sqrt;
  assign cyc_C3_sqrt = cyc_C3 & sqrtOp_PB;
  assign T222 = cyc_C6_sqrt | cyc_C5_div;
  assign cyc_C5_div = cyc_C5 & T223;
  assign T223 = sqrtOp_PB ^ 1'h1;
  assign cyc_C5 = T224;
  assign T224 = cycleNum_C == 3'h5;
  assign cyc_C6_sqrt = cycleNum_C == 3'h6;
  assign T225 = cyc_C4_sqrt | cyc_C2;
  assign cyc_C2 = T226;
  assign T226 = cycleNum_C == 3'h2;
  assign cyc_C4_sqrt = cyc_C4 & sqrtOp_PB;
  assign cyc_C4 = T227;
  assign T227 = cycleNum_C == 3'h4;
  assign T228 = T233 | T898;
  assign T898 = {1'h0, T229};
  assign T229 = cyc_C6_sqrt ? T230 : 104'h0;
  assign T230 = sigX1_B << 6'h2e;
  assign T231 = cyc_B3 ? sigXNU_B3_CX : sigX1_B;
  assign cyc_B3 = T232;
  assign T232 = cycleNum_B == 4'h3;
  assign T233 = cyc_B1 ? T234 : 105'h0;
  assign T234 = sigX1_B << 6'h2f;
  assign io_mulAddB_0 = T235;
  assign T235 = T899 | zComplSigT_C1;
  assign T899 = {1'h0, T236};
  assign T236 = T239 | T900;
  assign T900 = {20'h0, T237};
  assign T237 = cyc_C4 ? sqrSigma1_C : 33'h0;
  assign T238 = cyc_B1 ? sqrSigma1_B1 : sqrSigma1_C;
  assign sqrSigma1_B1 = io_mulAddResult_3[7'h4f:6'h2f];
  assign T239 = T242 | T901;
  assign T901 = {23'h0, T240};
  assign T240 = cyc_C6_sqrt ? T241 : 30'h0;
  assign T241 = sqrSigma1_C[5'h1e:1'h1];
  assign T242 = T246 | T902;
  assign T902 = {7'h0, zSigma1_B4};
  assign zSigma1_B4 = T243;
  assign T243 = cyc_B4 ? T244 : 46'h0;
  assign T244 = ~ T245;
  assign T245 = io_mulAddResult_3[7'h5a:6'h2d];
  assign T246 = T926 | T247;
  assign T247 = cyc_B6_sqrt ? T248 : 53'h0;
  assign T248 = ER1_B_sqrt << 6'h24;
  assign T249 = cyc_A1_sqrt ? ER1_A1_sqrt : ER1_B_sqrt;
  assign ER1_A1_sqrt = T467 ? T466 : T903;
  assign T903 = {1'h0, r1_A1};
  assign r1_A1 = {1'h1, fractR1_A1};
  assign fractR1_A1 = T250[4'he:1'h0];
  assign T250 = sqrtOp_PA ? T925 : T251;
  assign T251 = mulAdd9Out_A >> 4'h9;
  assign mulAdd9Out_A = {T460, T252};
  assign T252 = loMulAdd9Out_A[5'h11:1'h0];
  assign loMulAdd9Out_A = T917 + T253;
  assign T253 = {1'h0, T254};
  assign T254 = mulAdd9C_A[5'h11:1'h0];
  assign mulAdd9C_A = T271 | T904;
  assign T904 = {1'h0, T255};
  assign T255 = cyc_A1_div ? T256 : 24'h0;
  assign T256 = fractR0_A << 4'hf;
  assign T257 = T269 ? T258 : fractR0_A;
  assign T258 = zFractR0_A6_sqrt | zFractR0_A4_div;
  assign zFractR0_A4_div = T259[4'h8:1'h0];
  assign T259 = T262 ? T260 : 14'h0;
  assign T260 = T261 >> 4'hb;
  assign T261 = ~ mulAdd9Out_A;
  assign T262 = cyc_A4_div & T263;
  assign T263 = mulAdd9Out_A[5'h14];
  assign zFractR0_A6_sqrt = T264[4'h8:1'h0];
  assign T264 = T267 ? T265 : 15'h0;
  assign T265 = T266 >> 4'ha;
  assign T266 = ~ mulAdd9Out_A;
  assign T267 = cyc_A6_sqrt & T268;
  assign T268 = mulAdd9Out_A[5'h13];
  assign cyc_A6_sqrt = cycleNum_A == 3'h6;
  assign T269 = cyc_A6_sqrt | cyc_A4_div;
  assign cyc_A1_div = cyc_A1 & T270;
  assign T270 = sqrtOp_PA ^ 1'h1;
  assign T271 = T905 | T272;
  assign T272 = cyc_A1_sqrt ? T273 : 25'h0;
  assign T273 = fractR0_A << 5'h10;
  assign T905 = {4'h0, T274};
  assign T274 = T282 | T275;
  assign T275 = T281 ? partNegSigma0_A : 21'h0;
  assign T276 = T280 ? T277 : partNegSigma0_A;
  assign T277 = T278[5'h14:1'h0];
  assign T278 = cyc_A4_sqrt ? mulAdd9Out_A : T906;
  assign T906 = {9'h0, T279};
  assign T279 = mulAdd9Out_A >> 4'h9;
  assign cyc_A4_sqrt = cycleNum_A == 3'h4;
  assign T280 = cyc_A4_sqrt | cyc_A3;
  assign cyc_A3 = cycleNum_A == 3'h3;
  assign T281 = cyc_A3_sqrt | cyc_A2;
  assign cyc_A2 = cycleNum_A == 3'h2;
  assign cyc_A3_sqrt = cyc_A3 & sqrtOp_PA;
  assign T282 = T295 | T283;
  assign T283 = T287 ? T284 : 21'h0;
  assign T284 = T285 + 21'h400;
  assign T285 = sigB_PA[6'h2e:5'h1a];
  assign sigB_PA = {1'h1, T286};
  assign T286 = {fractB_51_PA, fractB_other_PA};
  assign T287 = T289 | cyc_A3_div;
  assign cyc_A3_div = cyc_A3 & T288;
  assign T288 = sqrtOp_PA ^ 1'h1;
  assign T289 = cyc_A4_sqrt & T290;
  assign T290 = hiSqrR0_A_sqrt[4'h9];
  assign T907 = T291[4'h9:1'h0];
  assign T291 = cyc_A5_sqrt ? T292 : T908;
  assign T908 = {6'h0, hiSqrR0_A_sqrt};
  assign T292 = sqrR0_A5_sqrt >> 4'ha;
  assign sqrR0_A5_sqrt = T294 ? T293 : T909;
  assign T909 = {1'h0, mulAdd9Out_A};
  assign T293 = mulAdd9Out_A << 1'h1;
  assign T294 = exp_PA[1'h0];
  assign cyc_A5_sqrt = cycleNum_A == 3'h5;
  assign T295 = T300 | T910;
  assign T910 = {10'h0, T296};
  assign T296 = T297 ? 11'h400 : 11'h0;
  assign T297 = cyc_A4_sqrt & T298;
  assign T298 = T299 ^ 1'h1;
  assign T299 = hiSqrR0_A_sqrt[4'h9];
  assign T300 = T304 | T911;
  assign T911 = {1'h0, T301};
  assign T301 = cyc_A5_sqrt ? T302 : 20'h0;
  assign T302 = 20'h40000 + T912;
  assign T912 = {1'h0, T303};
  assign T303 = fractR0_A << 4'ha;
  assign T304 = T914 | T305;
  assign T305 = {cyc_A4_div, T306};
  assign T306 = {zComplFractK0_A4_div, T307};
  assign T307 = 8'h0 - T913;
  assign T913 = {7'h0, cyc_A4_div};
  assign zComplFractK0_A4_div = T311 | T308;
  assign T308 = zLinPiece_7_A4_div ? 12'hef4 : 12'h0;
  assign zLinPiece_7_A4_div = cyc_A4_div & T309;
  assign T309 = T310 == 3'h7;
  assign T310 = fractB_S[6'h33:6'h31];
  assign T311 = T315 | T312;
  assign T312 = zLinPiece_6_A4_div ? 12'hdbd : 12'h0;
  assign zLinPiece_6_A4_div = cyc_A4_div & T313;
  assign T313 = T314 == 3'h6;
  assign T314 = fractB_S[6'h33:6'h31];
  assign T315 = T319 | T316;
  assign T316 = zLinPiece_5_A4_div ? 12'hc56 : 12'h0;
  assign zLinPiece_5_A4_div = cyc_A4_div & T317;
  assign T317 = T318 == 3'h5;
  assign T318 = fractB_S[6'h33:6'h31];
  assign T319 = T323 | T320;
  assign T320 = zLinPiece_4_A4_div ? 12'hab4 : 12'h0;
  assign zLinPiece_4_A4_div = cyc_A4_div & T321;
  assign T321 = T322 == 3'h4;
  assign T322 = fractB_S[6'h33:6'h31];
  assign T323 = T327 | T324;
  assign T324 = zLinPiece_3_A4_div ? 12'h8c6 : 12'h0;
  assign zLinPiece_3_A4_div = cyc_A4_div & T325;
  assign T325 = T326 == 3'h3;
  assign T326 = fractB_S[6'h33:6'h31];
  assign T327 = T331 | T328;
  assign T328 = zLinPiece_2_A4_div ? 12'h675 : 12'h0;
  assign zLinPiece_2_A4_div = cyc_A4_div & T329;
  assign T329 = T330 == 3'h2;
  assign T330 = fractB_S[6'h33:6'h31];
  assign T331 = T335 | T332;
  assign T332 = zLinPiece_1_A4_div ? 12'h3a2 : 12'h0;
  assign zLinPiece_1_A4_div = cyc_A4_div & T333;
  assign T333 = T334 == 3'h1;
  assign T334 = fractB_S[6'h33:6'h31];
  assign T335 = zLinPiece_0_A4_div ? 12'h1c : 12'h0;
  assign zLinPiece_0_A4_div = cyc_A4_div & T336;
  assign T336 = T337 == 3'h0;
  assign T337 = fractB_S[6'h33:6'h31];
  assign T914 = {1'h0, T338};
  assign T338 = T364 | T339;
  assign T339 = {cyc_A6_sqrt, T340};
  assign T340 = {zComplFractK0_A6_sqrt, T341};
  assign T341 = 6'h0 - T915;
  assign T915 = {5'h0, cyc_A6_sqrt};
  assign zComplFractK0_A6_sqrt = T346 | T342;
  assign T342 = zQuadPiece_3_A6_sqrt ? 13'h1b17 : 13'h0;
  assign zQuadPiece_3_A6_sqrt = T344 & T343;
  assign T343 = sigB_PA[6'h33];
  assign T344 = cyc_A6_sqrt & T345;
  assign T345 = exp_PA[1'h0];
  assign T346 = T352 | T347;
  assign T347 = zQuadPiece_2_A6_sqrt ? 13'h12d3 : 13'h0;
  assign zQuadPiece_2_A6_sqrt = T350 & T348;
  assign T348 = T349 ^ 1'h1;
  assign T349 = sigB_PA[6'h33];
  assign T350 = cyc_A6_sqrt & T351;
  assign T351 = exp_PA[1'h0];
  assign T352 = T358 | T353;
  assign T353 = zQuadPiece_1_A6_sqrt ? 13'hbca : 13'h0;
  assign zQuadPiece_1_A6_sqrt = T355 & T354;
  assign T354 = sigB_PA[6'h33];
  assign T355 = cyc_A6_sqrt & T356;
  assign T356 = T357 ^ 1'h1;
  assign T357 = exp_PA[1'h0];
  assign T358 = zQuadPiece_0_A6_sqrt ? 13'h1a : 13'h0;
  assign zQuadPiece_0_A6_sqrt = T361 & T359;
  assign T359 = T360 ^ 1'h1;
  assign T360 = sigB_PA[6'h33];
  assign T361 = cyc_A6_sqrt & T362;
  assign T362 = T363 ^ 1'h1;
  assign T363 = exp_PA[1'h0];
  assign T364 = {zComplK1_A7_sqrt, T365};
  assign T365 = 10'h0 - T916;
  assign T916 = {9'h0, cyc_A7_sqrt};
  assign zComplK1_A7_sqrt = T370 | T366;
  assign T366 = zQuadPiece_3_A7_sqrt ? 10'h27e : 10'h0;
  assign zQuadPiece_3_A7_sqrt = T368 & T367;
  assign T367 = fractB_S[6'h33];
  assign T368 = cyc_A7_sqrt & T369;
  assign T369 = expB_S[1'h0];
  assign T370 = T376 | T371;
  assign T371 = zQuadPiece_2_A7_sqrt ? 10'h14d : 10'h0;
  assign zQuadPiece_2_A7_sqrt = T374 & T372;
  assign T372 = T373 ^ 1'h1;
  assign T373 = fractB_S[6'h33];
  assign T374 = cyc_A7_sqrt & T375;
  assign T375 = expB_S[1'h0];
  assign T376 = T382 | T377;
  assign T377 = zQuadPiece_1_A7_sqrt ? 10'h1df : 10'h0;
  assign zQuadPiece_1_A7_sqrt = T379 & T378;
  assign T378 = fractB_S[6'h33];
  assign T379 = cyc_A7_sqrt & T380;
  assign T380 = T381 ^ 1'h1;
  assign T381 = expB_S[1'h0];
  assign T382 = zQuadPiece_0_A7_sqrt ? 10'h2f : 10'h0;
  assign zQuadPiece_0_A7_sqrt = T385 & T383;
  assign T383 = T384 ^ 1'h1;
  assign T384 = fractB_S[6'h33];
  assign T385 = cyc_A7_sqrt & T386;
  assign T386 = T387 ^ 1'h1;
  assign T387 = expB_S[1'h0];
  assign T917 = {1'h0, T388};
  assign T388 = mulAdd9A_A * mulAdd9B_A;
  assign mulAdd9B_A = T409 | T389;
  assign T389 = T408 ? nextMulAdd9B_A : 9'h0;
  assign T390 = T404 ? T391 : nextMulAdd9B_A;
  assign T391 = T395 | T392;
  assign T392 = cyc_A2 ? T393 : 9'h0;
  assign T393 = {1'h1, T394};
  assign T394 = fractR0_A[4'h8:1'h1];
  assign T395 = T398 | T396;
  assign T396 = cyc_A4_sqrt ? T397 : 9'h0;
  assign T397 = hiSqrR0_A_sqrt[4'h8:1'h0];
  assign T398 = T399 | zFractR0_A4_div;
  assign T399 = T402 | T400;
  assign T400 = cyc_A5_sqrt ? T401 : 9'h0;
  assign T401 = sqrR0_A5_sqrt[4'h9:1'h1];
  assign T402 = T403 | zFractR0_A6_sqrt;
  assign T403 = zFractB_A7_sqrt[6'h32:6'h2a];
  assign zFractB_A7_sqrt = cyc_A7_sqrt ? fractB_S : 52'h0;
  assign T404 = T405 | cyc_A2;
  assign T405 = T406 | cyc_A4;
  assign cyc_A4 = cyc_A4_sqrt | cyc_A4_div;
  assign T406 = T407 | cyc_A5_sqrt;
  assign T407 = cyc_A7_sqrt | cyc_A6_sqrt;
  assign T408 = cyc_S ^ 1'h1;
  assign T409 = zK1_A4_div | T410;
  assign T410 = zFractB_A7_sqrt[6'h32:6'h2a];
  assign zK1_A4_div = T412 | T411;
  assign T411 = zLinPiece_7_A4_div ? 9'h89 : 9'h0;
  assign T412 = T414 | T413;
  assign T413 = zLinPiece_6_A4_div ? 9'h9c : 9'h0;
  assign T414 = T416 | T415;
  assign T415 = zLinPiece_5_A4_div ? 9'hb4 : 9'h0;
  assign T416 = T418 | T417;
  assign T417 = zLinPiece_4_A4_div ? 9'hd2 : 9'h0;
  assign T418 = T420 | T419;
  assign T419 = zLinPiece_3_A4_div ? 9'hf8 : 9'h0;
  assign T420 = T422 | T421;
  assign T421 = zLinPiece_2_A4_div ? 9'h12a : 9'h0;
  assign T422 = T424 | T423;
  assign T423 = zLinPiece_1_A4_div ? 9'h16c : 9'h0;
  assign T424 = zLinPiece_0_A4_div ? 9'h1c7 : 9'h0;
  assign mulAdd9A_A = T452 | T425;
  assign T425 = T451 ? nextMulAdd9A_A : 9'h0;
  assign T918 = T426[4'h8:1'h0];
  assign T426 = T446 ? T427 : T919;
  assign T919 = {5'h0, nextMulAdd9A_A};
  assign T427 = T433 | T920;
  assign T920 = {5'h0, zSigma0_A2};
  assign zSigma0_A2 = T428[4'h8:1'h0];
  assign T428 = T431 ? T429 : 23'h0;
  assign T429 = T430 >> 2'h2;
  assign T430 = ~ mulAdd9Out_A;
  assign T431 = cyc_A2 & T432;
  assign T432 = mulAdd9Out_A[4'hb];
  assign T433 = T437 | T921;
  assign T921 = {5'h0, T434};
  assign T434 = T436 ? T435 : 9'h0;
  assign T435 = sigB_PA[6'h34:6'h2c];
  assign T436 = cyc_A5_sqrt | cyc_A3;
  assign T437 = T439 | T922;
  assign T922 = {5'h0, T438};
  assign T438 = zFractB_A4_div[6'h2b:6'h23];
  assign zFractB_A4_div = cyc_A4_div ? fractB_S : 52'h0;
  assign T439 = T442 | T923;
  assign T923 = {5'h0, T440};
  assign T440 = cyc_A4_sqrt ? T441 : 9'h0;
  assign T441 = sigB_PA[6'h2b:6'h23];
  assign T442 = T443 | T924;
  assign T924 = {5'h0, zFractR0_A6_sqrt};
  assign T443 = cyc_A7_sqrt ? T444 : 14'h0;
  assign T444 = T445 >> 4'hb;
  assign T445 = ~ mulAdd9Out_A;
  assign T446 = T447 | cyc_A2;
  assign T447 = T448 | cyc_A3;
  assign T448 = T449 | cyc_A4;
  assign T449 = T450 | cyc_A5_sqrt;
  assign T450 = cyc_A7_sqrt | cyc_A6_sqrt;
  assign T451 = cyc_S ^ 1'h1;
  assign T452 = T459 | zK2_A7_sqrt;
  assign zK2_A7_sqrt = T454 | T453;
  assign T453 = zQuadPiece_3_A7_sqrt ? 9'h89 : 9'h0;
  assign T454 = T456 | T455;
  assign T455 = zQuadPiece_2_A7_sqrt ? 9'h143 : 9'h0;
  assign T456 = T458 | T457;
  assign T457 = zQuadPiece_1_A7_sqrt ? 9'hc1 : 9'h0;
  assign T458 = zQuadPiece_0_A7_sqrt ? 9'h1c8 : 9'h0;
  assign T459 = zFractB_A4_div[6'h30:6'h28];
  assign T460 = T464 ? T462 : T461;
  assign T461 = mulAdd9C_A[5'h18:5'h12];
  assign T462 = T463 + 7'h1;
  assign T463 = mulAdd9C_A[5'h18:5'h12];
  assign T464 = loMulAdd9Out_A[5'h12];
  assign T925 = {1'h0, T465};
  assign T465 = mulAdd9Out_A >> 4'ha;
  assign T466 = r1_A1 << 1'h1;
  assign T467 = exp_PA[1'h0];
  assign cyc_A1_sqrt = cyc_A1 & sqrtOp_PA;
  assign cyc_B6_sqrt = T468;
  assign T468 = T469 & sqrtOp_PB;
  assign T469 = cyc_B6 & valid_PB;
  assign cyc_B6 = T470;
  assign T470 = cycleNum_B == 4'h6;
  assign T926 = {1'h0, T471};
  assign T471 = T476 | T927;
  assign T927 = {1'h0, T472};
  assign T472 = cyc_B7_sqrt ? T473 : 51'h0;
  assign T473 = ESqrR1_B_sqrt << 5'h13;
  assign T474 = cyc_B8_sqrt ? ESqrR1_B8_sqrt : ESqrR1_B_sqrt;
  assign ESqrR1_B8_sqrt = io_mulAddResult_3[7'h67:7'h48];
  assign cyc_B8_sqrt = T475;
  assign T475 = cycleNum_B == 4'h8;
  assign T476 = cyc_A1 ? T477 : 52'h0;
  assign T477 = r1_A1 << 6'h24;
  assign io_latchMulAddB_0 = T478;
  assign T478 = T479 | cyc_C1;
  assign T479 = T480 | cyc_C4;
  assign T480 = T481 | cyc_C6_sqrt;
  assign T481 = T482 | cyc_B4;
  assign T482 = T483 | cyc_B6_sqrt;
  assign T483 = cyc_A1 | cyc_B7_sqrt;
  assign io_mulAddA_0 = T484;
  assign T484 = T928 | zComplSigT_C1_sqrt;
  assign zComplSigT_C1_sqrt = T485;
  assign T485 = cyc_C1_sqrt ? T486 : 54'h0;
  assign T486 = ~ T487;
  assign T487 = io_mulAddResult_3[7'h68:6'h33];
  assign T928 = {1'h0, T488};
  assign T488 = T490 | T489;
  assign T489 = cyc_C1_div ? sigB_PC : 53'h0;
  assign T490 = T495 | T929;
  assign T929 = {7'h0, T491};
  assign T491 = cyc_C4_sqrt ? T492 : 46'h0;
  assign T492 = u_C_sqrt << 4'hf;
  assign T493 = cyc_C5_sqrt ? T494 : u_C_sqrt;
  assign T494 = sigXNU_B3_CX[6'h38:5'h1a];
  assign cyc_C5_sqrt = cyc_C5 & sqrtOp_PB;
  assign T495 = T500 | T930;
  assign T930 = {7'h0, T496};
  assign T496 = cyc_C4_div ? T497 : 46'h0;
  assign T497 = T498 << 4'hd;
  assign T498 = sigXN_C[6'h39:5'h19];
  assign cyc_C4_div = cyc_C4 & T499;
  assign T499 = sqrtOp_PB ^ 1'h1;
  assign T500 = T504 | T931;
  assign T931 = {7'h0, T501};
  assign T501 = T503 ? T502 : 46'h0;
  assign T502 = sigXNU_B3_CX[6'h39:4'hc];
  assign T503 = cyc_B3 | cyc_C6_sqrt;
  assign T504 = T506 | T932;
  assign T932 = {19'h0, T505};
  assign T505 = zSigma1_B4[6'h2d:4'hc];
  assign T506 = T514 | T507;
  assign T507 = cyc_B6_div ? sigA_PA : 53'h0;
  assign sigA_PA = {1'h1, T508};
  assign T508 = {fractA_51_PA, fractA_other_PA};
  assign T509 = T47 ? T510 : fractA_51_PA;
  assign T510 = fractA_S[6'h33];
  assign cyc_B6_div = T511;
  assign T511 = T513 & T512;
  assign T512 = sqrtOp_PA ^ 1'h1;
  assign T513 = cyc_B6 & valid_PA;
  assign T514 = T517 | T515;
  assign T515 = T516 ? sigB_PA : 53'h0;
  assign T516 = cyc_B7_sqrt | cyc_A1_div;
  assign T517 = cyc_A1_sqrt ? T518 : 53'h0;
  assign T518 = ER1_A1_sqrt << 6'h24;
  assign io_latchMulAddA_0 = T519;
  assign T519 = T520 | cyc_C1;
  assign T520 = T521 | cyc_C4;
  assign T521 = T522 | cyc_C6_sqrt;
  assign T522 = T523 | cyc_B3;
  assign T523 = T524 | cyc_B4;
  assign T524 = T525 | cyc_B6_div;
  assign T525 = cyc_A1 | cyc_B7_sqrt;
  assign io_usingMulAdd = T526;
  assign T526 = {T544, T527};
  assign T527 = {T532, T528};
  assign T528 = T531 | cyc_B2_sqrt;
  assign cyc_B2_sqrt = T529;
  assign T529 = cyc_B2 & sqrtOp_PB;
  assign cyc_B2 = T530;
  assign T530 = cycleNum_B == 4'h2;
  assign T531 = io_latchMulAddA_0 | cyc_B6;
  assign T532 = T533 | cyc_C2;
  assign T533 = T534 | cyc_C5;
  assign T534 = T536 | cyc_B1_sqrt;
  assign cyc_B1_sqrt = T535;
  assign T535 = cyc_B1 & sqrtOp_PB;
  assign T536 = T538 | cyc_B3_sqrt;
  assign cyc_B3_sqrt = T537;
  assign T537 = cyc_B3 & sqrtOp_PB;
  assign T538 = T539 | cyc_B4;
  assign T539 = T541 | cyc_B5;
  assign cyc_B5 = T540;
  assign T540 = cycleNum_B == 4'h5;
  assign T541 = T542 | cyc_B7_sqrt;
  assign T542 = T543 | cyc_B8_sqrt;
  assign T543 = cyc_A2 | cyc_A1_div;
  assign T544 = {T561, T545};
  assign T545 = T546 | cyc_C3;
  assign T546 = T547 | cyc_C6_sqrt;
  assign T547 = T550 | cyc_B1_div;
  assign cyc_B1_div = T548;
  assign T548 = cyc_B1 & T549;
  assign T549 = sqrtOp_PB ^ 1'h1;
  assign T550 = T551 | cyc_B2_sqrt;
  assign T551 = T554 | cyc_B4_sqrt;
  assign cyc_B4_sqrt = T552;
  assign T552 = T553 & sqrtOp_PB;
  assign T553 = cyc_B4 & valid_PB;
  assign T554 = T555 | cyc_B5;
  assign T555 = T556 | cyc_B6;
  assign T556 = T557 | cyc_B8_sqrt;
  assign T557 = T559 | cyc_B9_sqrt;
  assign cyc_B9_sqrt = T558;
  assign T558 = cycleNum_B == 4'h9;
  assign T559 = cyc_A3 | cyc_A2_div;
  assign cyc_A2_div = cyc_A2 & T560;
  assign T560 = sqrtOp_PA ^ 1'h1;
  assign T561 = T562 | cyc_C4;
  assign T562 = T563 | cyc_B1_sqrt;
  assign T563 = T566 | cyc_B2_div;
  assign cyc_B2_div = T564;
  assign T564 = cyc_B2 & T565;
  assign T565 = sqrtOp_PB ^ 1'h1;
  assign T566 = T567 | cyc_B3_sqrt;
  assign T567 = T570 | cyc_B5_sqrt;
  assign cyc_B5_sqrt = T568;
  assign T568 = T569 & sqrtOp_PB;
  assign T569 = cyc_B5 & valid_PB;
  assign T570 = T571 | cyc_B6;
  assign T571 = T572 | cyc_B7_sqrt;
  assign T572 = T573 | cyc_B9_sqrt;
  assign T573 = T575 | cyc_B10_sqrt;
  assign cyc_B10_sqrt = T574;
  assign T574 = cycleNum_B == 4'ha;
  assign T575 = T576 | cyc_A1_div;
  assign T576 = cyc_A4 | cyc_A3_div;
  assign io_exceptionFlags = T577;
  assign T577 = {T781, T578};
  assign T578 = {overflow_E1, T579};
  assign T579 = {underflow_E1, inexact_E1};
  assign inexact_E1 = T706 | T580;
  assign T580 = normalCase_PC & inexactY_E1;
  assign inexactY_E1 = hiRoundPosBit_E1 | anyRoundExtra_E1;
  assign anyRoundExtra_E1 = T677 | T581;
  assign T581 = all1sHiRoundExtraT_E ^ 1'h1;
  assign all1sHiRoundExtraT_E = T582 == 53'h0;
  assign T582 = T674 & T933;
  assign T933 = {1'h0, T583};
  assign T583 = roundMask_E >> 1'h1;
  assign roundMask_E = {T643, T584};
  assign T584 = {T618, T585};
  assign T585 = {T608, T586};
  assign T586 = T587[3'h4];
  assign T587 = T588[5'h14:5'h10];
  assign T588 = T589[6'h34:6'h20];
  assign T589 = T590[11'h402:10'h3ce];
  assign T590 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T591;
  assign T591 = ~ posExpX_E;
  assign posExpX_E = sExpX_E[4'hc:1'h0];
  assign sExpX_E = T595 | T934;
  assign T934 = {1'h0, T592};
  assign T592 = sqrtOp_PC ? T593 : 13'h0;
  assign T593 = T594 + 13'h400;
  assign T594 = exp_PC >> 1'h1;
  assign T595 = T605 | T596;
  assign T596 = T602 ? expP1_PC : 14'h0;
  assign expP1_PC = T601 ? T599 : T597;
  assign T597 = {T598, 1'h1};
  assign T598 = exp_PC[4'hd:1'h1];
  assign T599 = {T600, 1'h0};
  assign T600 = expP2_PC[4'hd:1'h1];
  assign expP2_PC = exp_PC + 14'h2;
  assign T601 = exp_PC[1'h0];
  assign T602 = T604 & T603;
  assign T603 = E_E_div ^ 1'h1;
  assign T604 = sqrtOp_PC ^ 1'h1;
  assign T605 = T606 ? exp_PC : 14'h0;
  assign T606 = T607 & E_E_div;
  assign T607 = sqrtOp_PC ^ 1'h1;
  assign T608 = {T614, T609};
  assign T609 = {T613, T610};
  assign T610 = T611[1'h1];
  assign T611 = T612[2'h3:2'h2];
  assign T612 = T587[2'h3:1'h0];
  assign T613 = T611[1'h0];
  assign T614 = {T617, T615};
  assign T615 = T616[1'h1];
  assign T616 = T612[1'h1:1'h0];
  assign T617 = T616[1'h0];
  assign T618 = T641 | T619;
  assign T619 = T620 & 16'haaaa;
  assign T620 = T621 << 1'h1;
  assign T621 = T622[4'he:1'h0];
  assign T622 = T639 | T623;
  assign T623 = T624 & 16'hcccc;
  assign T624 = T625 << 2'h2;
  assign T625 = T626[4'hd:1'h0];
  assign T626 = T637 | T627;
  assign T627 = T628 & 16'hf0f0;
  assign T628 = T629 << 3'h4;
  assign T629 = T630[4'hb:1'h0];
  assign T630 = T635 | T631;
  assign T631 = T632 & 16'hff00;
  assign T632 = T633 << 4'h8;
  assign T633 = T634[3'h7:1'h0];
  assign T634 = T588[4'hf:1'h0];
  assign T635 = T935 & 16'hff;
  assign T935 = {8'h0, T636};
  assign T636 = T634 >> 4'h8;
  assign T637 = T936 & 16'hf0f;
  assign T936 = {4'h0, T638};
  assign T638 = T630 >> 3'h4;
  assign T639 = T937 & 16'h3333;
  assign T937 = {2'h0, T640};
  assign T640 = T626 >> 2'h2;
  assign T641 = T938 & 16'h5555;
  assign T938 = {1'h0, T642};
  assign T642 = T622 >> 1'h1;
  assign T643 = T672 | T644;
  assign T644 = T645 & 32'haaaaaaaa;
  assign T645 = T646 << 1'h1;
  assign T646 = T647[5'h1e:1'h0];
  assign T647 = T670 | T648;
  assign T648 = T649 & 32'hcccccccc;
  assign T649 = T650 << 2'h2;
  assign T650 = T651[5'h1d:1'h0];
  assign T651 = T668 | T652;
  assign T652 = T653 & 32'hf0f0f0f0;
  assign T653 = T654 << 3'h4;
  assign T654 = T655[5'h1b:1'h0];
  assign T655 = T666 | T656;
  assign T656 = T657 & 32'hff00ff00;
  assign T657 = T658 << 4'h8;
  assign T658 = T659[5'h17:1'h0];
  assign T659 = T664 | T660;
  assign T660 = T661 & 32'hffff0000;
  assign T661 = T662 << 5'h10;
  assign T662 = T663[4'hf:1'h0];
  assign T663 = T589[5'h1f:1'h0];
  assign T664 = T939 & 32'hffff;
  assign T939 = {16'h0, T665};
  assign T665 = T663 >> 5'h10;
  assign T666 = T940 & 32'hff00ff;
  assign T940 = {8'h0, T667};
  assign T667 = T659 >> 4'h8;
  assign T668 = T941 & 32'hf0f0f0f;
  assign T941 = {4'h0, T669};
  assign T669 = T655 >> 3'h4;
  assign T670 = T942 & 32'h33333333;
  assign T942 = {2'h0, T671};
  assign T671 = T651 >> 2'h2;
  assign T672 = T943 & 32'h55555555;
  assign T943 = {1'h0, T673};
  assign T673 = T647 >> 1'h1;
  assign T674 = ~ sigT_E;
  assign T675 = cyc_C1 ? T676 : sigT_E;
  assign T676 = sigT_C1[6'h35:1'h1];
  assign T677 = T679 | T678;
  assign T678 = extraT_E ^ 1'h1;
  assign T679 = isZeroRemT_E ^ 1'h1;
  assign T680 = cyc_E2 ? T681 : isZeroRemT_E;
  assign T681 = T686 & T682;
  assign T682 = T685 | T683;
  assign T683 = T684 == 2'h0;
  assign T684 = remT_E2[6'h37:6'h36];
  assign remT_E2 = io_mulAddResult_3[6'h37:1'h0];
  assign T685 = sqrtOp_PC ^ 1'h1;
  assign T686 = T687 == 54'h0;
  assign T687 = remT_E2[6'h35:1'h0];
  assign cyc_E2 = T688;
  assign T688 = cycleNum_E == 3'h2;
  assign hiRoundPosBit_E1 = hiRoundPosBitT_E ^ T689;
  assign T689 = T690 & extraT_E;
  assign T690 = T691 & all1sHiRoundExtraT_E;
  assign T691 = T700 & T692;
  assign T692 = trueLtX_E1 ^ 1'h1;
  assign trueLtX_E1 = sqrtOp_PC ? T697 : isNegRemT_E;
  assign T693 = cyc_E2 ? T694 : isNegRemT_E;
  assign T694 = sqrtOp_PC ? T696 : T695;
  assign T695 = remT_E2[6'h35];
  assign T696 = remT_E2[6'h37];
  assign T697 = T699 & T698;
  assign T698 = isZeroRemT_E ^ 1'h1;
  assign T699 = isNegRemT_E ^ 1'h1;
  assign T700 = roundMask_E[1'h0];
  assign hiRoundPosBitT_E = T701 != 53'h0;
  assign T701 = sigT_E & T702;
  assign T702 = incrPosMask_E >> 1'h1;
  assign incrPosMask_E = T704 & T703;
  assign T703 = {roundMask_E, 1'h1};
  assign T704 = ~ T705;
  assign T705 = {1'h0, roundMask_E};
  assign T706 = overflow_E1 | underflow_E1;
  assign underflow_E1 = normalCase_PC & underflowY_E1;
  assign underflowY_E1 = totalUnderflowY_E1 | T707;
  assign T707 = T708 & inexactY_E1;
  assign T708 = posExpX_E <= 13'h401;
  assign totalUnderflowY_E1 = T776 | T709;
  assign T709 = T710 < 13'h3ce;
  assign T710 = sExpY_E1[4'hc:1'h0];
  assign sExpY_E1 = T760 | T944;
  assign T944 = {1'h0, T711};
  assign T711 = T714 ? T712 : 13'h0;
  assign T712 = T713 + 13'h400;
  assign T713 = expP2_PC >> 1'h1;
  assign T714 = T715 & sqrtOp_PC;
  assign T715 = sigY_E1[6'h35];
  assign sigY_E1 = T725 & T716;
  assign T716 = ~ roundEvenMask_E1;
  assign roundEvenMask_E1 = T717 ? incrPosMask_E : 54'h0;
  assign T717 = T719 & T718;
  assign T718 = anyRoundExtra_E1 ^ 1'h1;
  assign T719 = roundingMode_near_even_PC & hiRoundPosBit_E1;
  assign roundingMode_near_even_PC = roundingMode_PC == 2'h0;
  assign T720 = entering_PC ? T721 : roundingMode_PC;
  assign T721 = valid_PB ? roundingMode_PB : io_roundingMode;
  assign T722 = entering_PB ? T723 : roundingMode_PB;
  assign T723 = valid_PA ? roundingMode_PA : io_roundingMode;
  assign T724 = entering_PA ? io_roundingMode : roundingMode_PA;
  assign T725 = T731 ? sigY1_E : sigY0_E;
  assign sigY0_E = sigAdjT_E & T726;
  assign T726 = {1'h1, T727};
  assign T727 = ~ roundMask_E;
  assign sigAdjT_E = T728 + T945;
  assign T945 = {53'h0, roundMagUp_PC};
  assign roundMagUp_PC = sign_PC ? roundingMode_min_PC : roundingMode_max_PC;
  assign roundingMode_max_PC = roundingMode_PC == 2'h3;
  assign roundingMode_min_PC = roundingMode_PC == 2'h2;
  assign T728 = 54'h0 + T946;
  assign T946 = {1'h0, sigT_E};
  assign sigY1_E = T729 + 54'h1;
  assign T729 = sigAdjT_E | T730;
  assign T730 = {1'h0, roundMask_E};
  assign T731 = T743 | T732;
  assign T732 = roundingMode_near_even_PC & T733;
  assign T733 = T737 | T734;
  assign T734 = T735 & all1sHiRoundExtraT_E;
  assign T735 = extraT_E & T736;
  assign T736 = trueLtX_E1 ^ 1'h1;
  assign T737 = hiRoundPosBitT_E | T738;
  assign T738 = T741 & T739;
  assign T739 = T740 ^ 1'h1;
  assign T740 = roundMask_E[1'h0];
  assign T741 = extraT_E | T742;
  assign T742 = trueLtX_E1 ^ 1'h1;
  assign T743 = T754 | T744;
  assign T744 = roundMagUp_PC & T745;
  assign T745 = T750 | T746;
  assign T746 = all1sHiRoundT_E ^ 1'h1;
  assign all1sHiRoundT_E = T747 & all1sHiRoundExtraT_E;
  assign T747 = T748 | hiRoundPosBitT_E;
  assign T748 = T749 ^ 1'h1;
  assign T749 = roundMask_E[1'h0];
  assign T750 = T752 & T751;
  assign T751 = isZeroRemT_E ^ 1'h1;
  assign T752 = extraT_E & T753;
  assign T753 = trueLtX_E1 ^ 1'h1;
  assign T754 = T755 & all1sHiRoundT_E;
  assign T755 = T757 & T756;
  assign T756 = trueLtX_E1 ^ 1'h1;
  assign T757 = roundMagDown_PC & extraT_E;
  assign roundMagDown_PC = T759 & T758;
  assign T758 = roundingMode_near_even_PC ^ 1'h1;
  assign T759 = roundMagUp_PC ^ 1'h1;
  assign T760 = T767 | T761;
  assign T761 = T762 ? expP2_PC : 14'h0;
  assign T762 = T764 & T763;
  assign T763 = E_E_div ^ 1'h1;
  assign T764 = T766 & T765;
  assign T765 = sqrtOp_PC ^ 1'h1;
  assign T766 = sigY_E1[6'h35];
  assign T767 = T773 | T768;
  assign T768 = T769 ? expP1_PC : 14'h0;
  assign T769 = T770 & E_E_div;
  assign T770 = T772 & T771;
  assign T771 = sqrtOp_PC ^ 1'h1;
  assign T772 = sigY_E1[6'h35];
  assign T773 = T774 ? sExpX_E : 14'h0;
  assign T774 = T775 ^ 1'h1;
  assign T775 = sigY_E1[6'h35];
  assign T776 = sExpY_E1[4'hd];
  assign overflow_E1 = normalCase_PC & overflowY_E1;
  assign overflowY_E1 = T779 & T777;
  assign T777 = 3'h3 <= T778;
  assign T778 = sExpY_E1[4'hc:4'ha];
  assign T779 = T780 ^ 1'h1;
  assign T780 = sExpY_E1[4'hd];
  assign T781 = {invalid_PC, infinity_PC};
  assign infinity_PC = T782 & isZeroB_PC;
  assign T782 = T784 & T783;
  assign T783 = isZeroA_PC ^ 1'h1;
  assign T784 = T786 & T785;
  assign T785 = isSpecialA_PC ^ 1'h1;
  assign T786 = sqrtOp_PC ^ 1'h1;
  assign invalid_PC = T799 | notSigNaN_invalid_PC;
  assign notSigNaN_invalid_PC = sqrtOp_PC ? T794 : T787;
  assign T787 = T793 | T788;
  assign T788 = isInfA_PC & isInfB_PC;
  assign isInfB_PC = isSpecialB_PC & T789;
  assign T789 = T790 ^ 1'h1;
  assign T790 = specialCodeB_PC[1'h0];
  assign isInfA_PC = isSpecialA_PC & T791;
  assign T791 = T792 ^ 1'h1;
  assign T792 = specialCodeA_PC[1'h0];
  assign T793 = isZeroA_PC & isZeroB_PC;
  assign T794 = T795 & sign_PC;
  assign T795 = T797 & T796;
  assign T796 = isZeroB_PC ^ 1'h1;
  assign T797 = isNaNB_PC ^ 1'h1;
  assign isNaNB_PC = isSpecialB_PC & T798;
  assign T798 = specialCodeB_PC[1'h0];
  assign T799 = T801 | isSigNaNB_PC;
  assign isSigNaNB_PC = isNaNB_PC & T800;
  assign T800 = fractB_51_PC ^ 1'h1;
  assign T801 = T810 & isSigNaNA_PC;
  assign isSigNaNA_PC = isNaNA_PC & T802;
  assign T802 = fractA_51_PC ^ 1'h1;
  assign T803 = entering_PC ? T804 : fractA_51_PC;
  assign T804 = valid_PB ? fractA_51_PB : T805;
  assign T805 = fractA_S[6'h33];
  assign T806 = entering_PB ? T807 : fractA_51_PB;
  assign T807 = valid_PA ? fractA_51_PA : T808;
  assign T808 = fractA_S[6'h33];
  assign isNaNA_PC = isSpecialA_PC & T809;
  assign T809 = specialCodeA_PC[1'h0];
  assign T810 = sqrtOp_PC ^ 1'h1;
  assign io_out = T811;
  assign T811 = {signOut_PC, T812};
  assign T812 = {expOut_E1, fractOut_E1};
  assign fractOut_E1 = T815 | T813;
  assign T813 = 52'h0 - T947;
  assign T947 = {51'h0, pegMaxFiniteMagOut_E1};
  assign pegMaxFiniteMagOut_E1 = overflow_E1 & T814;
  assign T814 = overflowY_roundMagUp_PC ^ 1'h1;
  assign overflowY_roundMagUp_PC = roundingMode_near_even_PC | roundMagUp_PC;
  assign T815 = T820 ? T816 : fractY_E1;
  assign fractY_E1 = sigY_E1[6'h33:1'h0];
  assign T816 = isNaNOut_PC ? 52'h8000000000000 : 52'h0;
  assign isNaNOut_PC = T817 | notSigNaN_invalid_PC;
  assign T817 = T818 | isNaNB_PC;
  assign T818 = T819 & isNaNA_PC;
  assign T819 = sqrtOp_PC ^ 1'h1;
  assign T820 = T821 | isNaNOut_PC;
  assign T821 = notSpecial_isZeroOut_E1 | totalUnderflowY_E1;
  assign notSpecial_isZeroOut_E1 = sqrtOp_PC ? isZeroB_PC : T822;
  assign T822 = T825 | T823;
  assign T823 = totalUnderflowY_E1 & T824;
  assign T824 = roundMagUp_PC ^ 1'h1;
  assign T825 = isZeroA_PC | isInfB_PC;
  assign expOut_E1 = T827 | T826;
  assign T826 = isNaNOut_PC ? 12'he00 : 12'h0;
  assign T827 = T832 | T828;
  assign T828 = notNaN_isInfOut_E1 ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut_E1 = sqrtOp_PC ? isInfB_PC : T829;
  assign T829 = T831 | T830;
  assign T830 = overflow_E1 & overflowY_roundMagUp_PC;
  assign T831 = isInfA_PC | isZeroB_PC;
  assign T832 = T834 | T833;
  assign T833 = pegMaxFiniteMagOut_E1 ? 12'hbff : 12'h0;
  assign T834 = T837 | T835;
  assign T835 = pegMinFiniteMagOut_E1 ? 12'h3ce : 12'h0;
  assign pegMinFiniteMagOut_E1 = T836 & roundMagUp_PC;
  assign T836 = normalCase_PC & totalUnderflowY_E1;
  assign T837 = T840 & T838;
  assign T838 = ~ T839;
  assign T839 = notNaN_isInfOut_E1 ? 12'h200 : 12'h0;
  assign T840 = T843 & T841;
  assign T841 = ~ T842;
  assign T842 = pegMaxFiniteMagOut_E1 ? 12'h400 : 12'h0;
  assign T843 = T846 & T844;
  assign T844 = ~ T845;
  assign T845 = pegMinFiniteMagOut_E1 ? 12'hc31 : 12'h0;
  assign T846 = expY_E1 & T847;
  assign T847 = ~ T848;
  assign T848 = notSpecial_isZeroOut_E1 ? 12'he00 : 12'h0;
  assign expY_E1 = sExpY_E1[4'hb:1'h0];
  assign signOut_PC = T851 & T849;
  assign T849 = sqrtOp_PC ? T850 : sign_PC;
  assign T850 = isZeroB_PC & sign_PC;
  assign T851 = isNaNOut_PC ^ 1'h1;
  assign io_outValid_sqrt = T852;
  assign T852 = leaving_PC & sqrtOp_PC;
  assign io_outValid_div = T853;
  assign T853 = leaving_PC & T854;
  assign T854 = sqrtOp_PC ^ 1'h1;
  assign io_inReady_sqrt = T855;
  assign T855 = T857 & T856;
  assign T856 = cyc_B1_sqrt ^ 1'h1;
  assign T857 = T859 & T858;
  assign T858 = cyc_B2_div ^ 1'h1;
  assign T859 = T861 & T860;
  assign T860 = cyc_B4_sqrt ^ 1'h1;
  assign T861 = T863 & T862;
  assign T862 = cyc_B5_sqrt ^ 1'h1;
  assign T863 = ready_PA & T864;
  assign T864 = cyc_B6_sqrt ^ 1'h1;
  assign ready_PA = T865;
  assign T865 = T866 | valid_leaving_PA;
  assign T866 = valid_PA ^ 1'h1;
  assign io_inReady_div = T867;
  assign T867 = T869 & T868;
  assign T868 = cyc_C4 ^ 1'h1;
  assign T869 = T871 & T870;
  assign T870 = cyc_C5 ^ 1'h1;
  assign T871 = T873 & T872;
  assign T872 = cyc_B1_sqrt ^ 1'h1;
  assign T873 = T875 & T874;
  assign T874 = cyc_B2 ^ 1'h1;
  assign T875 = T877 & T876;
  assign T876 = cyc_B3 ^ 1'h1;
  assign T877 = T879 & T878;
  assign T878 = cyc_B4_sqrt ^ 1'h1;
  assign T879 = T881 & T880;
  assign T880 = cyc_B5_sqrt ^ 1'h1;
  assign T881 = T883 & T882;
  assign T882 = cyc_B6_sqrt ^ 1'h1;
  assign T883 = ready_PA & T884;
  assign T884 = cyc_B7_sqrt ^ 1'h1;

  always @(posedge clk) begin
    if(cyc_C1) begin
      extraT_E <= T7;
    end
    if(entering_PC) begin
      sqrtOp_PC <= T17;
    end
    if(entering_PB) begin
      sqrtOp_PB <= T19;
    end
    if(entering_PA) begin
      sqrtOp_PA <= io_sqrtOp;
    end
    if(reset) begin
      cycleNum_E <= 3'h0;
    end else if(T30) begin
      cycleNum_E <= T28;
    end
    if(entering_PC) begin
      specialCodeB_PC <= T36;
    end
    if(entering_PB) begin
      specialCodeB_PB <= T38;
    end
    if(entering_PA) begin
      specialCodeB_PA <= specialCodeB_S;
    end
    if(entering_PC) begin
      specialCodeA_PC <= T43;
    end
    if(entering_PB) begin
      specialCodeA_PB <= T45;
    end
    if(T47) begin
      specialCodeA_PA <= specialCodeA_S;
    end
    if(entering_PC) begin
      sign_PC <= T57;
    end
    if(entering_PB) begin
      sign_PB <= T60;
    end
    if(entering_PA) begin
      sign_PA <= sign_S;
    end
    if(reset) begin
      valid_PC <= 1'h0;
    end else if(T67) begin
      valid_PC <= entering_PC;
    end
    if(reset) begin
      cycleNum_C <= 3'h0;
    end else if(T106) begin
      cycleNum_C <= T71;
    end
    if(reset) begin
      cycleNum_B <= 4'h0;
    end else if(T104) begin
      cycleNum_B <= T76;
    end
    if(reset) begin
      cycleNum_A <= 3'h0;
    end else if(T102) begin
      cycleNum_A <= T80;
    end
    if(reset) begin
      valid_PA <= 1'h0;
    end else if(T124) begin
      valid_PA <= entering_PA;
    end
    if(reset) begin
      valid_PB <= 1'h0;
    end else if(T155) begin
      valid_PB <= entering_PB;
    end
    if(entering_PC_normalCase) begin
      fractB_other_PC <= fractB_other_PB;
    end
    if(entering_PB_normalCase) begin
      fractB_other_PB <= fractB_other_PA;
    end
    if(entering_PA_normalCase) begin
      fractB_other_PA <= T176;
    end
    if(entering_PC) begin
      fractB_51_PC <= T180;
    end
    if(entering_PB) begin
      fractB_51_PB <= T183;
    end
    if(entering_PA) begin
      fractB_51_PA <= T186;
    end
    if(entering_PC_normalCase) begin
      exp_PC <= exp_PB;
    end
    if(entering_PB_normalCase) begin
      exp_PB <= exp_PA;
    end
    if(entering_PA_normalCase) begin
      exp_PA <= T196;
    end
    if(entering_PC_normalCase) begin
      fractA_0_PC <= fractA_0_PB;
    end
    if(entering_PB_normalCase) begin
      fractA_0_PB <= T209;
    end
    if(cyc_A4_div) begin
      fractA_other_PA <= T211;
    end
    if(cyc_C1) begin
      E_E_div <= E_C1_div;
    end
    if(T221) begin
      sigXN_C <= sigXNU_B3_CX;
    end
    if(cyc_B3) begin
      sigX1_B <= sigXNU_B3_CX;
    end
    if(cyc_B1) begin
      sqrSigma1_C <= sqrSigma1_B1;
    end
    if(cyc_A1_sqrt) begin
      ER1_B_sqrt <= ER1_A1_sqrt;
    end
    if(T269) begin
      fractR0_A <= T258;
    end
    if(T280) begin
      partNegSigma0_A <= T277;
    end
    hiSqrR0_A_sqrt <= T907;
    if(T404) begin
      nextMulAdd9B_A <= T391;
    end
    nextMulAdd9A_A <= T918;
    if(cyc_B8_sqrt) begin
      ESqrR1_B_sqrt <= ESqrR1_B8_sqrt;
    end
    if(cyc_C5_sqrt) begin
      u_C_sqrt <= T494;
    end
    if(T47) begin
      fractA_51_PA <= T510;
    end
    if(cyc_C1) begin
      sigT_E <= T676;
    end
    if(cyc_E2) begin
      isZeroRemT_E <= T681;
    end
    if(cyc_E2) begin
      isNegRemT_E <= T694;
    end
    if(entering_PC) begin
      roundingMode_PC <= T721;
    end
    if(entering_PB) begin
      roundingMode_PB <= T723;
    end
    if(entering_PA) begin
      roundingMode_PA <= io_roundingMode;
    end
    if(entering_PC) begin
      fractA_51_PC <= T804;
    end
    if(entering_PB) begin
      fractA_51_PB <= T807;
    end
  end
endmodule

module Mul54(input clk,
    input  io_val_s0,
    input  io_latch_a_s0,
    input [53:0] io_a_s0,
    input  io_latch_b_s0,
    input [53:0] io_b_s0,
    input [104:0] io_c_s2,
    output[104:0] io_result_s3
);

  reg [104:0] reg_result_s3;
  wire[104:0] T0;
  wire[104:0] T1;
  wire[104:0] T2;
  wire[107:0] T3;
  reg [53:0] reg_b_s2;
  wire[53:0] T4;
  reg [53:0] reg_b_s1;
  wire[53:0] T5;
  wire T6;
  reg  val_s1;
  reg [53:0] reg_a_s2;
  wire[53:0] T7;
  reg [53:0] reg_a_s1;
  wire[53:0] T8;
  wire T9;
  reg  val_s2;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_result_s3 = {4{$random}};
    reg_b_s2 = {2{$random}};
    reg_b_s1 = {2{$random}};
    val_s1 = {1{$random}};
    reg_a_s2 = {2{$random}};
    reg_a_s1 = {2{$random}};
    val_s2 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_result_s3 = reg_result_s3;
  assign T0 = val_s2 ? T1 : reg_result_s3;
  assign T1 = T2 + io_c_s2;
  assign T2 = T3[7'h68:1'h0];
  assign T3 = reg_a_s2 * reg_b_s2;
  assign T4 = val_s1 ? reg_b_s1 : reg_b_s2;
  assign T5 = T6 ? io_b_s0 : reg_b_s1;
  assign T6 = io_val_s0 & io_latch_b_s0;
  assign T7 = val_s1 ? reg_a_s1 : reg_a_s2;
  assign T8 = T9 ? io_a_s0 : reg_a_s1;
  assign T9 = io_val_s0 & io_latch_a_s0;

  always @(posedge clk) begin
    if(val_s2) begin
      reg_result_s3 <= T1;
    end
    if(val_s1) begin
      reg_b_s2 <= reg_b_s1;
    end
    if(T6) begin
      reg_b_s1 <= io_b_s0;
    end
    val_s1 <= io_val_s0;
    if(val_s1) begin
      reg_a_s2 <= reg_a_s1;
    end
    if(T9) begin
      reg_a_s1 <= io_a_s0;
    end
    val_s2 <= val_s1;
  end
endmodule

module DivSqrtRecF64(input clk, input reset,
    output io_inReady_div,
    output io_inReady_sqrt,
    input  io_inValid,
    input  io_sqrtOp,
    input [64:0] io_a,
    input [64:0] io_b,
    input [1:0] io_roundingMode,
    output io_outValid_div,
    output io_outValid_sqrt,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire T0;
  wire ds_io_inReady_div;
  wire ds_io_inReady_sqrt;
  wire ds_io_outValid_div;
  wire ds_io_outValid_sqrt;
  wire[64:0] ds_io_out;
  wire[4:0] ds_io_exceptionFlags;
  wire[3:0] ds_io_usingMulAdd;
  wire ds_io_latchMulAddA_0;
  wire[53:0] ds_io_mulAddA_0;
  wire ds_io_latchMulAddB_0;
  wire[53:0] ds_io_mulAddB_0;
  wire[104:0] ds_io_mulAddC_2;
  wire[104:0] mul_io_result_s3;


  assign T0 = ds_io_usingMulAdd[1'h0];
  assign io_exceptionFlags = ds_io_exceptionFlags;
  assign io_out = ds_io_out;
  assign io_outValid_sqrt = ds_io_outValid_sqrt;
  assign io_outValid_div = ds_io_outValid_div;
  assign io_inReady_sqrt = ds_io_inReady_sqrt;
  assign io_inReady_div = ds_io_inReady_div;
  DivSqrtRecF64_mulAddZ31 ds(.clk(clk), .reset(reset),
       .io_inReady_div( ds_io_inReady_div ),
       .io_inReady_sqrt( ds_io_inReady_sqrt ),
       .io_inValid( io_inValid ),
       .io_sqrtOp( io_sqrtOp ),
       .io_a( io_a ),
       .io_b( io_b ),
       .io_roundingMode( io_roundingMode ),
       .io_outValid_div( ds_io_outValid_div ),
       .io_outValid_sqrt( ds_io_outValid_sqrt ),
       .io_out( ds_io_out ),
       .io_exceptionFlags( ds_io_exceptionFlags ),
       .io_usingMulAdd( ds_io_usingMulAdd ),
       .io_latchMulAddA_0( ds_io_latchMulAddA_0 ),
       .io_mulAddA_0( ds_io_mulAddA_0 ),
       .io_latchMulAddB_0( ds_io_latchMulAddB_0 ),
       .io_mulAddB_0( ds_io_mulAddB_0 ),
       .io_mulAddC_2( ds_io_mulAddC_2 ),
       .io_mulAddResult_3( mul_io_result_s3 )
  );
  Mul54 mul(.clk(clk),
       .io_val_s0( T0 ),
       .io_latch_a_s0( ds_io_latchMulAddA_0 ),
       .io_a_s0( ds_io_mulAddA_0 ),
       .io_latch_b_s0( ds_io_latchMulAddB_0 ),
       .io_b_s0( ds_io_mulAddB_0 ),
       .io_c_s2( ds_io_mulAddC_2 ),
       .io_result_s3( mul_io_result_s3 )
  );
endmodule

module FPU(input clk, input reset,
    input [31:0] io_inst,
    input [63:0] io_fromint_data,
    input [2:0] io_fcsr_rm,
    output io_fcsr_flags_valid,
    output[4:0] io_fcsr_flags_bits,
    output[63:0] io_store_data,
    output[63:0] io_toint_data,
    input  io_dmem_resp_val,
    input [2:0] io_dmem_resp_type,
    input [4:0] io_dmem_resp_tag,
    input [63:0] io_dmem_resp_data,
    input  io_valid,
    output io_fcsr_rdy,
    output io_nack_mem,
    output io_illegal_rm,
    input  io_killx,
    input  io_killm,
    output[4:0] io_dec_cmd,
    output io_dec_ldst,
    output io_dec_wen,
    output io_dec_ren1,
    output io_dec_ren2,
    output io_dec_ren3,
    output io_dec_swap12,
    output io_dec_swap23,
    output io_dec_single,
    output io_dec_fromint,
    output io_dec_toint,
    output io_dec_fastpipe,
    output io_dec_fma,
    output io_dec_div,
    output io_dec_sqrt,
    output io_dec_round,
    output io_dec_wflags,
    output io_sboard_set,
    output io_sboard_clr,
    output[4:0] io_sboard_clra,
    output io_cp_req_ready,
    input  io_cp_req_valid,
    input [4:0] io_cp_req_bits_cmd,
    input  io_cp_req_bits_ldst,
    input  io_cp_req_bits_wen,
    input  io_cp_req_bits_ren1,
    input  io_cp_req_bits_ren2,
    input  io_cp_req_bits_ren3,
    input  io_cp_req_bits_swap12,
    input  io_cp_req_bits_swap23,
    input  io_cp_req_bits_single,
    input  io_cp_req_bits_fromint,
    input  io_cp_req_bits_toint,
    input  io_cp_req_bits_fastpipe,
    input  io_cp_req_bits_fma,
    input  io_cp_req_bits_div,
    input  io_cp_req_bits_sqrt,
    input  io_cp_req_bits_round,
    input  io_cp_req_bits_wflags,
    input [2:0] io_cp_req_bits_rm,
    input [1:0] io_cp_req_bits_typ,
    input [64:0] io_cp_req_bits_in1,
    input [64:0] io_cp_req_bits_in2,
    input [64:0] io_cp_req_bits_in3,
    input  io_cp_resp_ready,
    output io_cp_resp_valid,
    output[64:0] io_cp_resp_bits_data
    //output[4:0] io_cp_resp_bits_exc
);

  reg [1:0] R0;
  wire[1:0] T1;
  wire T2;
  wire divSqrt_inReady;
  wire T3;
  reg [64:0] R4;
  wire[64:0] T5;
  wire T6;
  wire[1:0] T339;
  reg  mem_ctrl_sqrt;
  wire T7;
  wire T8;
  wire cp_ctrl_sqrt;
  reg  R9;
  wire T10;
  reg  ex_reg_valid;
  wire T340;
  wire req_valid;
  wire T11;
  wire T12;
  reg  divSqrt_in_flight;
  wire T341;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg  mem_ctrl_div;
  wire T17;
  wire T18;
  wire cp_ctrl_div;
  reg  R19;
  wire T20;
  reg  mem_reg_valid;
  wire T342;
  wire T21;
  wire ex_cp_valid;
  wire T22;
  wire T23;
  wire T24;
  wire[64:0] req_in3;
  wire[64:0] T25;
  wire[64:0] cp_rs3;
  wire[64:0] ex_rs3;
  reg [64:0] regfile [31:0];
  wire[64:0] T26;
  wire[64:0] wdata;
  wire[64:0] T27;
  wire[64:0] T28;
  wire T29;
  wire[1:0] T30;
  wire[1:0] T343;
  wire[2:0] wsrc;
  reg [8:0] winfo_0;
  wire[8:0] T31;
  wire[8:0] T32;
  reg [8:0] winfo_1;
  wire[8:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] memLatencyMask;
  wire[1:0] T37;
  wire T38;
  wire T39;
  reg  mem_ctrl_single;
  wire T40;
  wire T41;
  wire cp_ctrl_single;
  reg  R42;
  wire T43;
  reg  mem_ctrl_fma;
  wire T44;
  wire T45;
  wire cp_ctrl_fma;
  reg  R46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T344;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  reg  mem_ctrl_fromint;
  wire T52;
  wire T53;
  wire cp_ctrl_fromint;
  reg  R54;
  wire T55;
  wire[1:0] T345;
  reg  mem_ctrl_fastpipe;
  wire T56;
  wire T57;
  wire cp_ctrl_fastpipe;
  reg  R58;
  wire T59;
  wire T60;
  reg  write_port_busy;
  wire T61;
  wire T62;
  wire T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] T66;
  wire T67;
  wire T68;
  wire[3:0] T69;
  wire[3:0] T346;
  wire[2:0] T70;
  wire T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[3:0] T347;
  wire[2:0] T74;
  wire[3:0] T348;
  reg [1:0] wen;
  wire[1:0] T349;
  wire[1:0] T75;
  wire[1:0] T350;
  wire T76;
  wire[1:0] T77;
  wire[1:0] T351;
  wire T78;
  wire T79;
  wire T80;
  wire killm;
  wire T81;
  reg  mem_cp_valid;
  wire T352;
  wire T82;
  wire T83;
  wire T84;
  wire[2:0] T85;
  wire[2:0] T86;
  wire[2:0] T87;
  wire T88;
  wire T89;
  wire[2:0] T90;
  wire[2:0] T353;
  wire[1:0] T91;
  wire T92;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T354;
  wire[1:0] T95;
  wire[2:0] T355;
  wire mem_wen;
  wire T96;
  wire T97;
  wire T98;
  wire[8:0] mem_winfo;
  wire[5:0] T99;
  wire[4:0] T100;
  reg [31:0] mem_reg_inst;
  wire[31:0] T101;
  reg [31:0] ex_reg_inst;
  wire[31:0] T102;
  wire[2:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire T110;
  wire[1:0] T356;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[64:0] T116;
  wire T117;
  wire T118;
  wire[64:0] divSqrt_wdata;
  wire[64:0] T119;
  wire[64:0] T357;
  reg  R120;
  wire T121;
  reg  divSqrt_wen;
  wire T122;
  wire T123;
  reg  divSqrt_killed;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire wcp;
  wire[4:0] waddr;
  wire[4:0] T129;
  wire[4:0] T130;
  reg [4:0] divSqrt_waddr;
  wire[4:0] T131;
  wire[4:0] T132;
  wire[64:0] T133;
  wire[64:0] load_wb_data_recoded;
  wire[64:0] rec_d;
  wire[63:0] T134;
  wire[51:0] T135;
  wire[51:0] T136;
  reg [63:0] load_wb_data;
  wire[63:0] T137;
  wire[51:0] T138;
  wire[50:0] T139;
  wire[114:0] T140;
  wire[5:0] T141;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[5:0] T365;
  wire[5:0] T366;
  wire[5:0] T367;
  wire[5:0] T368;
  wire[5:0] T369;
  wire[5:0] T370;
  wire[5:0] T371;
  wire[5:0] T372;
  wire[5:0] T373;
  wire[5:0] T374;
  wire[5:0] T375;
  wire[5:0] T376;
  wire[5:0] T377;
  wire[5:0] T378;
  wire[5:0] T379;
  wire[5:0] T380;
  wire[5:0] T381;
  wire[5:0] T382;
  wire[5:0] T383;
  wire[5:0] T384;
  wire[5:0] T385;
  wire[5:0] T386;
  wire[5:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[4:0] T392;
  wire[4:0] T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire[4:0] T396;
  wire[4:0] T397;
  wire[4:0] T398;
  wire[4:0] T399;
  wire[4:0] T400;
  wire[4:0] T401;
  wire[4:0] T402;
  wire[4:0] T403;
  wire[4:0] T404;
  wire[4:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire[3:0] T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[2:0] T414;
  wire[2:0] T415;
  wire[2:0] T416;
  wire[2:0] T417;
  wire[1:0] T418;
  wire[1:0] T419;
  wire T420;
  wire[63:0] T143;
  wire[63:0] T144;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T145;
  wire[10:0] T146;
  wire[11:0] T147;
  wire[11:0] T483;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  wire[11:0] T154;
  wire[11:0] T484;
  wire[10:0] T155;
  wire[10:0] T485;
  wire[1:0] T156;
  wire[11:0] T157;
  wire[11:0] T486;
  wire[11:0] T158;
  wire[11:0] T487;
  wire[11:0] T159;
  wire[11:0] T160;
  wire[11:0] T161;
  wire[2:0] T162;
  wire[2:0] T488;
  wire T163;
  wire T164;
  wire[64:0] T165;
  wire[32:0] rec_s;
  wire[31:0] T166;
  wire[22:0] T167;
  wire[22:0] T168;
  wire[22:0] T169;
  wire[21:0] T170;
  wire[53:0] T171;
  wire[4:0] T172;
  wire[4:0] T489;
  wire[4:0] T490;
  wire[4:0] T491;
  wire[4:0] T492;
  wire[4:0] T493;
  wire[4:0] T494;
  wire[4:0] T495;
  wire[4:0] T496;
  wire[4:0] T497;
  wire[4:0] T498;
  wire[4:0] T499;
  wire[4:0] T500;
  wire[4:0] T501;
  wire[4:0] T502;
  wire[4:0] T503;
  wire[4:0] T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[3:0] T510;
  wire[3:0] T511;
  wire[3:0] T512;
  wire[2:0] T513;
  wire[2:0] T514;
  wire[2:0] T515;
  wire[2:0] T516;
  wire[1:0] T517;
  wire[1:0] T518;
  wire T519;
  wire[31:0] T174;
  wire[31:0] T175;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T176;
  wire[7:0] T177;
  wire[8:0] T178;
  wire[8:0] T550;
  wire[6:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[8:0] T185;
  wire[8:0] T551;
  wire[7:0] T186;
  wire[7:0] T552;
  wire[1:0] T187;
  wire[8:0] T188;
  wire[8:0] T553;
  wire[8:0] T189;
  wire[8:0] T554;
  wire[8:0] T190;
  wire[8:0] T191;
  wire[8:0] T192;
  wire[2:0] T193;
  wire[2:0] T555;
  wire T194;
  wire T195;
  reg  load_wb_single;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg  load_wb;
  reg [4:0] load_wb_tag;
  wire[4:0] T200;
  reg [4:0] ex_ra3;
  wire[4:0] T201;
  wire[4:0] T202;
  wire[4:0] T203;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire[64:0] req_in2;
  wire[64:0] T208;
  wire[64:0] cp_rs2;
  wire[64:0] ex_rs2;
  reg [4:0] ex_ra2;
  wire[4:0] T209;
  wire[4:0] T210;
  wire[4:0] T211;
  wire T212;
  wire T213;
  wire[4:0] T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire[64:0] req_in1;
  wire[64:0] T219;
  wire[64:0] ex_rs1;
  reg [4:0] ex_ra1;
  wire[4:0] T220;
  wire[4:0] T221;
  wire[4:0] T222;
  wire T223;
  wire T224;
  wire[4:0] T225;
  wire T226;
  wire[1:0] req_typ;
  wire[1:0] T227;
  wire[1:0] T228;
  wire[2:0] req_rm;
  wire[2:0] T229;
  wire[2:0] ex_rm;
  wire[2:0] T230;
  wire T231;
  wire[2:0] T232;
  wire req_wflags;
  wire T233;
  wire cp_ctrl_wflags;
  reg  R234;
  wire T235;
  wire req_round;
  wire T236;
  wire cp_ctrl_round;
  reg  R237;
  wire T238;
  wire req_sqrt;
  wire req_div;
  wire req_fma;
  wire req_fastpipe;
  wire req_toint;
  wire T239;
  wire cp_ctrl_toint;
  reg  R240;
  wire T241;
  wire req_fromint;
  wire req_single;
  wire req_swap23;
  wire T242;
  wire cp_ctrl_swap23;
  reg  R243;
  wire T244;
  wire req_swap12;
  wire T245;
  wire cp_ctrl_swap12;
  reg  R246;
  wire T247;
  wire req_ren3;
  wire T248;
  wire cp_ctrl_ren3;
  reg  R249;
  wire T250;
  wire req_ren2;
  wire T251;
  wire cp_ctrl_ren2;
  reg  R252;
  wire T253;
  wire req_ren1;
  wire T254;
  wire cp_ctrl_ren1;
  reg  R255;
  wire T256;
  wire req_wen;
  wire T257;
  wire cp_ctrl_wen;
  reg  R258;
  wire T259;
  wire req_ldst;
  wire T260;
  wire cp_ctrl_ldst;
  reg  R261;
  wire T262;
  wire[4:0] req_cmd;
  wire[4:0] T263;
  wire[4:0] cp_ctrl_cmd;
  reg [4:0] R264;
  wire[4:0] T265;
  wire T266;
  wire[64:0] T267;
  wire[64:0] T556;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[64:0] T280;
  wire[64:0] T557;
  wire[63:0] T281;
  wire T282;
  reg  mem_ctrl_toint;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  reg  wb_cp_valid;
  wire T558;
  wire T291;
  reg  R292;
  wire T293;
  wire T294;
  wire T295;
  reg  wb_reg_valid;
  wire T559;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire units_busy;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  reg  wb_ctrl_toint;
  wire T314;
  wire T315;
  wire T316;
  reg  mem_ctrl_wflags;
  wire T317;
  wire T318;
  wire[4:0] T319;
  wire[4:0] T320;
  wire[4:0] wexc;
  wire[4:0] T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T560;
  wire[4:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire[4:0] T328;
  wire[4:0] T329;
  wire[4:0] divSqrt_flags;
  wire[4:0] T330;
  wire[4:0] T331;
  reg [4:0] R332;
  wire[4:0] T333;
  wire[4:0] T334;
  reg [4:0] wb_toint_exc;
  wire[4:0] T335;
  wire wb_toint_valid;
  wire T336;
  wire T337;
  wire T338;
  wire[4:0] fp_decoder_io_sigs_cmd;
  wire fp_decoder_io_sigs_ldst;
  wire fp_decoder_io_sigs_wen;
  wire fp_decoder_io_sigs_ren1;
  wire fp_decoder_io_sigs_ren2;
  wire fp_decoder_io_sigs_ren3;
  wire fp_decoder_io_sigs_swap12;
  wire fp_decoder_io_sigs_swap23;
  wire fp_decoder_io_sigs_single;
  wire fp_decoder_io_sigs_fromint;
  wire fp_decoder_io_sigs_toint;
  wire fp_decoder_io_sigs_fastpipe;
  wire fp_decoder_io_sigs_fma;
  wire fp_decoder_io_sigs_div;
  wire fp_decoder_io_sigs_sqrt;
  wire fp_decoder_io_sigs_round;
  wire fp_decoder_io_sigs_wflags;
  wire[2:0] fpiu_io_as_double_rm;
  wire[64:0] fpiu_io_as_double_in1;
  wire[64:0] fpiu_io_as_double_in2;
  wire fpiu_io_out_valid;
  wire fpiu_io_out_bits_lt;
  wire[63:0] fpiu_io_out_bits_store;
  wire[63:0] fpiu_io_out_bits_toint;
  wire[4:0] fpiu_io_out_bits_exc;
  wire[64:0] ifpu_io_out_bits_data;
  wire[4:0] ifpu_io_out_bits_exc;
  wire DivSqrtRecF64_io_inReady_div;
  wire DivSqrtRecF64_io_inReady_sqrt;
  wire DivSqrtRecF64_io_outValid_div;
  wire DivSqrtRecF64_io_outValid_sqrt;
  wire[64:0] DivSqrtRecF64_io_out;
  wire[4:0] DivSqrtRecF64_io_exceptionFlags;
  wire[32:0] RecFNToRecFN_io_out;
  wire[4:0] RecFNToRecFN_io_exceptionFlags;
  wire[64:0] sfma_io_out_bits_data;
  wire[4:0] sfma_io_out_bits_exc;
  wire[64:0] dfma_io_out_bits_data;
  wire[4:0] dfma_io_out_bits_exc;
  wire[64:0] fpmu_io_out_bits_data;
  wire[4:0] fpmu_io_out_bits_exc;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R4 = {3{$random}};
    mem_ctrl_sqrt = {1{$random}};
    R9 = {1{$random}};
    ex_reg_valid = {1{$random}};
    divSqrt_in_flight = {1{$random}};
    mem_ctrl_div = {1{$random}};
    R19 = {1{$random}};
    mem_reg_valid = {1{$random}};
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      regfile[initvar] = {3{$random}};
    winfo_0 = {1{$random}};
    winfo_1 = {1{$random}};
    mem_ctrl_single = {1{$random}};
    R42 = {1{$random}};
    mem_ctrl_fma = {1{$random}};
    R46 = {1{$random}};
    mem_ctrl_fromint = {1{$random}};
    R54 = {1{$random}};
    mem_ctrl_fastpipe = {1{$random}};
    R58 = {1{$random}};
    write_port_busy = {1{$random}};
    wen = {1{$random}};
    mem_cp_valid = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    R120 = {1{$random}};
    divSqrt_wen = {1{$random}};
    divSqrt_killed = {1{$random}};
    divSqrt_waddr = {1{$random}};
    load_wb_data = {2{$random}};
    load_wb_single = {1{$random}};
    load_wb = {1{$random}};
    load_wb_tag = {1{$random}};
    ex_ra3 = {1{$random}};
    ex_ra2 = {1{$random}};
    ex_ra1 = {1{$random}};
    R234 = {1{$random}};
    R237 = {1{$random}};
    R240 = {1{$random}};
    R243 = {1{$random}};
    R246 = {1{$random}};
    R249 = {1{$random}};
    R252 = {1{$random}};
    R255 = {1{$random}};
    R258 = {1{$random}};
    R261 = {1{$random}};
    R264 = {1{$random}};
    mem_ctrl_toint = {1{$random}};
    wb_cp_valid = {1{$random}};
    R292 = {1{$random}};
    wb_reg_valid = {1{$random}};
    wb_ctrl_toint = {1{$random}};
    mem_ctrl_wflags = {1{$random}};
    R332 = {1{$random}};
    wb_toint_exc = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_cp_resp_bits_exc = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 ? T339 : R0;
  assign T2 = T11 & divSqrt_inReady;
  assign divSqrt_inReady = T3;
  assign T3 = mem_ctrl_sqrt ? DivSqrtRecF64_io_inReady_sqrt : DivSqrtRecF64_io_inReady_div;
  assign T5 = T6 ? DivSqrtRecF64_io_out : R4;
  assign T6 = DivSqrtRecF64_io_outValid_div | DivSqrtRecF64_io_outValid_sqrt;
  assign T339 = fpiu_io_as_double_rm[1'h1:1'h0];
  assign T7 = req_valid ? T8 : mem_ctrl_sqrt;
  assign T8 = ex_reg_valid ? R9 : cp_ctrl_sqrt;
  assign cp_ctrl_sqrt = io_cp_req_bits_sqrt;
  assign T10 = io_valid ? fp_decoder_io_sigs_sqrt : R9;
  assign T340 = reset ? 1'h0 : io_valid;
  assign req_valid = ex_reg_valid | io_cp_req_valid;
  assign T11 = T15 & T12;
  assign T12 = divSqrt_in_flight ^ 1'h1;
  assign T341 = reset ? 1'h0 : T13;
  assign T13 = T6 ? 1'h0 : T14;
  assign T14 = T2 ? 1'h1 : divSqrt_in_flight;
  assign T15 = mem_reg_valid & T16;
  assign T16 = mem_ctrl_div | mem_ctrl_sqrt;
  assign T17 = req_valid ? T18 : mem_ctrl_div;
  assign T18 = ex_reg_valid ? R19 : cp_ctrl_div;
  assign cp_ctrl_div = io_cp_req_bits_div;
  assign T20 = io_valid ? fp_decoder_io_sigs_div : R19;
  assign T342 = reset ? 1'h0 : T21;
  assign T21 = T23 | ex_cp_valid;
  assign ex_cp_valid = io_cp_req_valid & T22;
  assign T22 = ex_reg_valid ^ 1'h1;
  assign T23 = ex_reg_valid & T24;
  assign T24 = io_killx ^ 1'h1;
  assign req_in3 = T25;
  assign T25 = ex_reg_valid ? ex_rs3 : cp_rs3;
  assign cp_rs3 = io_cp_req_bits_swap23 ? io_cp_req_bits_in2 : io_cp_req_bits_in3;
  assign ex_rs3 = regfile[ex_ra3];
  assign wdata = divSqrt_wen ? divSqrt_wdata : T27;
  assign T27 = T118 ? T116 : T28;
  assign T28 = T29 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T29 = T30[1'h0];
  assign T30 = T343;
  assign T343 = wsrc[1'h1:1'h0];
  assign wsrc = winfo_0 >> 3'h6;
  assign T31 = T112 ? mem_winfo : T32;
  assign T32 = T98 ? winfo_1 : winfo_0;
  assign T33 = T34 ? mem_winfo : winfo_1;
  assign T34 = mem_wen & T35;
  assign T35 = T60 & T36;
  assign T36 = memLatencyMask[1'h1];
  assign memLatencyMask = T48 | T37;
  assign T37 = T38 ? 2'h2 : 2'h0;
  assign T38 = mem_ctrl_fma & T39;
  assign T39 = mem_ctrl_single ^ 1'h1;
  assign T40 = req_valid ? T41 : mem_ctrl_single;
  assign T41 = ex_reg_valid ? R42 : cp_ctrl_single;
  assign cp_ctrl_single = io_cp_req_bits_single;
  assign T43 = io_valid ? fp_decoder_io_sigs_single : R42;
  assign T44 = req_valid ? T45 : mem_ctrl_fma;
  assign T45 = ex_reg_valid ? R46 : cp_ctrl_fma;
  assign cp_ctrl_fma = io_cp_req_bits_fma;
  assign T47 = io_valid ? fp_decoder_io_sigs_fma : R46;
  assign T48 = T50 | T344;
  assign T344 = {1'h0, T49};
  assign T49 = mem_ctrl_fma & mem_ctrl_single;
  assign T50 = T345 | T51;
  assign T51 = mem_ctrl_fromint ? 2'h2 : 2'h0;
  assign T52 = req_valid ? T53 : mem_ctrl_fromint;
  assign T53 = ex_reg_valid ? R54 : cp_ctrl_fromint;
  assign cp_ctrl_fromint = io_cp_req_bits_fromint;
  assign T55 = io_valid ? fp_decoder_io_sigs_fromint : R54;
  assign T345 = {1'h0, mem_ctrl_fastpipe};
  assign T56 = req_valid ? T57 : mem_ctrl_fastpipe;
  assign T57 = ex_reg_valid ? R58 : cp_ctrl_fastpipe;
  assign cp_ctrl_fastpipe = io_cp_req_bits_fastpipe;
  assign T59 = io_valid ? fp_decoder_io_sigs_fastpipe : R58;
  assign T60 = write_port_busy ^ 1'h1;
  assign T61 = req_valid ? T62 : write_port_busy;
  assign T62 = T83 | T63;
  assign T63 = T64 != 4'h0;
  assign T64 = T348 & T65;
  assign T65 = T69 | T66;
  assign T66 = T67 ? 4'h8 : 4'h0;
  assign T67 = T45 & T68;
  assign T68 = T41 ^ 1'h1;
  assign T69 = T72 | T346;
  assign T346 = {1'h0, T70};
  assign T70 = T71 ? 3'h4 : 3'h0;
  assign T71 = T45 & T41;
  assign T72 = T347 | T73;
  assign T73 = T53 ? 4'h8 : 4'h0;
  assign T347 = {1'h0, T74};
  assign T74 = T57 ? 3'h4 : 3'h0;
  assign T348 = {2'h0, wen};
  assign T349 = reset ? 2'h0 : T75;
  assign T75 = T79 ? T77 : T350;
  assign T350 = {1'h0, T76};
  assign T76 = wen >> 1'h1;
  assign T77 = T351 | memLatencyMask;
  assign T351 = {1'h0, T78};
  assign T78 = wen >> 1'h1;
  assign T79 = mem_wen & T80;
  assign T80 = killm ^ 1'h1;
  assign killm = T82 & T81;
  assign T81 = mem_cp_valid ^ 1'h1;
  assign T352 = reset ? 1'h0 : ex_cp_valid;
  assign T82 = io_killm | io_nack_mem;
  assign T83 = mem_wen & T84;
  assign T84 = T85 != 3'h0;
  assign T85 = T355 & T86;
  assign T86 = T90 | T87;
  assign T87 = T88 ? 3'h4 : 3'h0;
  assign T88 = T45 & T89;
  assign T89 = T41 ^ 1'h1;
  assign T90 = T93 | T353;
  assign T353 = {1'h0, T91};
  assign T91 = T92 ? 2'h2 : 2'h0;
  assign T92 = T45 & T41;
  assign T93 = T354 | T94;
  assign T94 = T53 ? 3'h4 : 3'h0;
  assign T354 = {1'h0, T95};
  assign T95 = T57 ? 2'h2 : 2'h0;
  assign T355 = {1'h0, memLatencyMask};
  assign mem_wen = mem_reg_valid & T96;
  assign T96 = T97 | mem_ctrl_fromint;
  assign T97 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T98 = wen[1'h1];
  assign mem_winfo = {T103, T99};
  assign T99 = {mem_ctrl_single, T100};
  assign T100 = mem_reg_inst[4'hb:3'h7];
  assign T101 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T102 = io_valid ? io_inst : ex_reg_inst;
  assign T103 = {mem_cp_valid, T104};
  assign T104 = T108 | T105;
  assign T105 = T106 ? 2'h3 : 2'h0;
  assign T106 = mem_ctrl_fma & T107;
  assign T107 = mem_ctrl_single ^ 1'h1;
  assign T108 = T356 | T109;
  assign T109 = T110 ? 2'h2 : 2'h0;
  assign T110 = mem_ctrl_fma & mem_ctrl_single;
  assign T356 = {1'h0, T111};
  assign T111 = 1'h0 | mem_ctrl_fromint;
  assign T112 = mem_wen & T113;
  assign T113 = T115 & T114;
  assign T114 = memLatencyMask[1'h0];
  assign T115 = write_port_busy ^ 1'h1;
  assign T116 = T117 ? dfma_io_out_bits_data : sfma_io_out_bits_data;
  assign T117 = T30[1'h0];
  assign T118 = T30[1'h1];
  assign divSqrt_wdata = T119;
  assign T119 = R120 ? T357 : R4;
  assign T357 = {32'h0, RecFNToRecFN_io_out};
  assign T121 = T2 ? mem_ctrl_single : R120;
  assign T122 = T6 ? T123 : 1'h0;
  assign T123 = divSqrt_killed ^ 1'h1;
  assign T124 = T2 ? killm : divSqrt_killed;
  assign T125 = T126 | divSqrt_wen;
  assign T126 = T128 & T127;
  assign T127 = wen[1'h0];
  assign T128 = wcp ^ 1'h1;
  assign wcp = winfo_0[4'h8];
  assign waddr = divSqrt_wen ? divSqrt_waddr : T129;
  assign T129 = T130;
  assign T130 = winfo_0[3'h4:1'h0];
  assign T131 = T2 ? T132 : divSqrt_waddr;
  assign T132 = mem_reg_inst[4'hb:3'h7];
  assign load_wb_data_recoded = load_wb_single ? T165 : rec_d;
  assign rec_d = {T164, T134};
  assign T134 = {T147, T135};
  assign T135 = T145 ? T138 : T136;
  assign T136 = load_wb_data[6'h33:1'h0];
  assign T137 = io_dmem_resp_val ? io_dmem_resp_data : load_wb_data;
  assign T138 = {T139, 1'h0};
  assign T139 = T140[6'h32:1'h0];
  assign T140 = T136 << T141;
  assign T141 = ~ T358;
  assign T358 = T482 ? 6'h3f : T359;
  assign T359 = T481 ? 6'h3e : T360;
  assign T360 = T480 ? 6'h3d : T361;
  assign T361 = T479 ? 6'h3c : T362;
  assign T362 = T478 ? 6'h3b : T363;
  assign T363 = T477 ? 6'h3a : T364;
  assign T364 = T476 ? 6'h39 : T365;
  assign T365 = T475 ? 6'h38 : T366;
  assign T366 = T474 ? 6'h37 : T367;
  assign T367 = T473 ? 6'h36 : T368;
  assign T368 = T472 ? 6'h35 : T369;
  assign T369 = T471 ? 6'h34 : T370;
  assign T370 = T470 ? 6'h33 : T371;
  assign T371 = T469 ? 6'h32 : T372;
  assign T372 = T468 ? 6'h31 : T373;
  assign T373 = T467 ? 6'h30 : T374;
  assign T374 = T466 ? 6'h2f : T375;
  assign T375 = T465 ? 6'h2e : T376;
  assign T376 = T464 ? 6'h2d : T377;
  assign T377 = T463 ? 6'h2c : T378;
  assign T378 = T462 ? 6'h2b : T379;
  assign T379 = T461 ? 6'h2a : T380;
  assign T380 = T460 ? 6'h29 : T381;
  assign T381 = T459 ? 6'h28 : T382;
  assign T382 = T458 ? 6'h27 : T383;
  assign T383 = T457 ? 6'h26 : T384;
  assign T384 = T456 ? 6'h25 : T385;
  assign T385 = T455 ? 6'h24 : T386;
  assign T386 = T454 ? 6'h23 : T387;
  assign T387 = T453 ? 6'h22 : T388;
  assign T388 = T452 ? 6'h21 : T389;
  assign T389 = T451 ? 6'h20 : T390;
  assign T390 = T450 ? 5'h1f : T391;
  assign T391 = T449 ? 5'h1e : T392;
  assign T392 = T448 ? 5'h1d : T393;
  assign T393 = T447 ? 5'h1c : T394;
  assign T394 = T446 ? 5'h1b : T395;
  assign T395 = T445 ? 5'h1a : T396;
  assign T396 = T444 ? 5'h19 : T397;
  assign T397 = T443 ? 5'h18 : T398;
  assign T398 = T442 ? 5'h17 : T399;
  assign T399 = T441 ? 5'h16 : T400;
  assign T400 = T440 ? 5'h15 : T401;
  assign T401 = T439 ? 5'h14 : T402;
  assign T402 = T438 ? 5'h13 : T403;
  assign T403 = T437 ? 5'h12 : T404;
  assign T404 = T436 ? 5'h11 : T405;
  assign T405 = T435 ? 5'h10 : T406;
  assign T406 = T434 ? 4'hf : T407;
  assign T407 = T433 ? 4'he : T408;
  assign T408 = T432 ? 4'hd : T409;
  assign T409 = T431 ? 4'hc : T410;
  assign T410 = T430 ? 4'hb : T411;
  assign T411 = T429 ? 4'ha : T412;
  assign T412 = T428 ? 4'h9 : T413;
  assign T413 = T427 ? 4'h8 : T414;
  assign T414 = T426 ? 3'h7 : T415;
  assign T415 = T425 ? 3'h6 : T416;
  assign T416 = T424 ? 3'h5 : T417;
  assign T417 = T423 ? 3'h4 : T418;
  assign T418 = T422 ? 2'h3 : T419;
  assign T419 = T421 ? 2'h2 : T420;
  assign T420 = T143[1'h1];
  assign T143 = T144;
  assign T144 = T136 << 4'hc;
  assign T421 = T143[2'h2];
  assign T422 = T143[2'h3];
  assign T423 = T143[3'h4];
  assign T424 = T143[3'h5];
  assign T425 = T143[3'h6];
  assign T426 = T143[3'h7];
  assign T427 = T143[4'h8];
  assign T428 = T143[4'h9];
  assign T429 = T143[4'ha];
  assign T430 = T143[4'hb];
  assign T431 = T143[4'hc];
  assign T432 = T143[4'hd];
  assign T433 = T143[4'he];
  assign T434 = T143[4'hf];
  assign T435 = T143[5'h10];
  assign T436 = T143[5'h11];
  assign T437 = T143[5'h12];
  assign T438 = T143[5'h13];
  assign T439 = T143[5'h14];
  assign T440 = T143[5'h15];
  assign T441 = T143[5'h16];
  assign T442 = T143[5'h17];
  assign T443 = T143[5'h18];
  assign T444 = T143[5'h19];
  assign T445 = T143[5'h1a];
  assign T446 = T143[5'h1b];
  assign T447 = T143[5'h1c];
  assign T448 = T143[5'h1d];
  assign T449 = T143[5'h1e];
  assign T450 = T143[5'h1f];
  assign T451 = T143[6'h20];
  assign T452 = T143[6'h21];
  assign T453 = T143[6'h22];
  assign T454 = T143[6'h23];
  assign T455 = T143[6'h24];
  assign T456 = T143[6'h25];
  assign T457 = T143[6'h26];
  assign T458 = T143[6'h27];
  assign T459 = T143[6'h28];
  assign T460 = T143[6'h29];
  assign T461 = T143[6'h2a];
  assign T462 = T143[6'h2b];
  assign T463 = T143[6'h2c];
  assign T464 = T143[6'h2d];
  assign T465 = T143[6'h2e];
  assign T466 = T143[6'h2f];
  assign T467 = T143[6'h30];
  assign T468 = T143[6'h31];
  assign T469 = T143[6'h32];
  assign T470 = T143[6'h33];
  assign T471 = T143[6'h34];
  assign T472 = T143[6'h35];
  assign T473 = T143[6'h36];
  assign T474 = T143[6'h37];
  assign T475 = T143[6'h38];
  assign T476 = T143[6'h39];
  assign T477 = T143[6'h3a];
  assign T478 = T143[6'h3b];
  assign T479 = T143[6'h3c];
  assign T480 = T143[6'h3d];
  assign T481 = T143[6'h3e];
  assign T482 = T143[6'h3f];
  assign T145 = T146 == 11'h0;
  assign T146 = load_wb_data[6'h3e:6'h34];
  assign T147 = T159 | T483;
  assign T483 = {2'h0, T148};
  assign T148 = T149 << 4'h9;
  assign T149 = T152 & T150;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T136 == 52'h0;
  assign T152 = T153 == 2'h3;
  assign T153 = T154[4'hb:4'ha];
  assign T154 = T157 + T484;
  assign T484 = {1'h0, T155};
  assign T155 = 11'h400 | T485;
  assign T485 = {9'h0, T156};
  assign T156 = T145 ? 2'h2 : 2'h1;
  assign T157 = T145 ? T158 : T486;
  assign T486 = {1'h0, T146};
  assign T158 = T487 ^ 12'hfff;
  assign T487 = {6'h0, T141};
  assign T159 = T154 & T160;
  assign T160 = ~ T161;
  assign T161 = T162 << 4'h9;
  assign T162 = 3'h0 - T488;
  assign T488 = {2'h0, T163};
  assign T163 = T145 & T151;
  assign T164 = load_wb_data[6'h3f];
  assign T165 = {32'hffffffff, rec_s};
  assign rec_s = {T195, T166};
  assign T166 = {T178, T167};
  assign T167 = T176 ? T169 : T168;
  assign T168 = load_wb_data[5'h16:1'h0];
  assign T169 = {T170, 1'h0};
  assign T170 = T171[5'h15:1'h0];
  assign T171 = T168 << T172;
  assign T172 = ~ T489;
  assign T489 = T549 ? 5'h1f : T490;
  assign T490 = T548 ? 5'h1e : T491;
  assign T491 = T547 ? 5'h1d : T492;
  assign T492 = T546 ? 5'h1c : T493;
  assign T493 = T545 ? 5'h1b : T494;
  assign T494 = T544 ? 5'h1a : T495;
  assign T495 = T543 ? 5'h19 : T496;
  assign T496 = T542 ? 5'h18 : T497;
  assign T497 = T541 ? 5'h17 : T498;
  assign T498 = T540 ? 5'h16 : T499;
  assign T499 = T539 ? 5'h15 : T500;
  assign T500 = T538 ? 5'h14 : T501;
  assign T501 = T537 ? 5'h13 : T502;
  assign T502 = T536 ? 5'h12 : T503;
  assign T503 = T535 ? 5'h11 : T504;
  assign T504 = T534 ? 5'h10 : T505;
  assign T505 = T533 ? 4'hf : T506;
  assign T506 = T532 ? 4'he : T507;
  assign T507 = T531 ? 4'hd : T508;
  assign T508 = T530 ? 4'hc : T509;
  assign T509 = T529 ? 4'hb : T510;
  assign T510 = T528 ? 4'ha : T511;
  assign T511 = T527 ? 4'h9 : T512;
  assign T512 = T526 ? 4'h8 : T513;
  assign T513 = T525 ? 3'h7 : T514;
  assign T514 = T524 ? 3'h6 : T515;
  assign T515 = T523 ? 3'h5 : T516;
  assign T516 = T522 ? 3'h4 : T517;
  assign T517 = T521 ? 2'h3 : T518;
  assign T518 = T520 ? 2'h2 : T519;
  assign T519 = T174[1'h1];
  assign T174 = T175;
  assign T175 = T168 << 4'h9;
  assign T520 = T174[2'h2];
  assign T521 = T174[2'h3];
  assign T522 = T174[3'h4];
  assign T523 = T174[3'h5];
  assign T524 = T174[3'h6];
  assign T525 = T174[3'h7];
  assign T526 = T174[4'h8];
  assign T527 = T174[4'h9];
  assign T528 = T174[4'ha];
  assign T529 = T174[4'hb];
  assign T530 = T174[4'hc];
  assign T531 = T174[4'hd];
  assign T532 = T174[4'he];
  assign T533 = T174[4'hf];
  assign T534 = T174[5'h10];
  assign T535 = T174[5'h11];
  assign T536 = T174[5'h12];
  assign T537 = T174[5'h13];
  assign T538 = T174[5'h14];
  assign T539 = T174[5'h15];
  assign T540 = T174[5'h16];
  assign T541 = T174[5'h17];
  assign T542 = T174[5'h18];
  assign T543 = T174[5'h19];
  assign T544 = T174[5'h1a];
  assign T545 = T174[5'h1b];
  assign T546 = T174[5'h1c];
  assign T547 = T174[5'h1d];
  assign T548 = T174[5'h1e];
  assign T549 = T174[5'h1f];
  assign T176 = T177 == 8'h0;
  assign T177 = load_wb_data[5'h1e:5'h17];
  assign T178 = T190 | T550;
  assign T550 = {2'h0, T179};
  assign T179 = T180 << 3'h6;
  assign T180 = T183 & T181;
  assign T181 = T182 ^ 1'h1;
  assign T182 = T168 == 23'h0;
  assign T183 = T184 == 2'h3;
  assign T184 = T185[4'h8:3'h7];
  assign T185 = T188 + T551;
  assign T551 = {1'h0, T186};
  assign T186 = 8'h80 | T552;
  assign T552 = {6'h0, T187};
  assign T187 = T176 ? 2'h2 : 2'h1;
  assign T188 = T176 ? T189 : T553;
  assign T553 = {1'h0, T177};
  assign T189 = T554 ^ 9'h1ff;
  assign T554 = {4'h0, T172};
  assign T190 = T185 & T191;
  assign T191 = ~ T192;
  assign T192 = T193 << 3'h6;
  assign T193 = 3'h0 - T555;
  assign T555 = {2'h0, T194};
  assign T194 = T176 & T182;
  assign T195 = load_wb_data[5'h1f];
  assign T196 = io_dmem_resp_val ? T197 : load_wb_single;
  assign T197 = T199 | T198;
  assign T198 = io_dmem_resp_type == 3'h6;
  assign T199 = io_dmem_resp_type == 3'h2;
  assign T200 = io_dmem_resp_val ? io_dmem_resp_tag : load_wb_tag;
  assign T201 = T207 ? T206 : T202;
  assign T202 = T204 ? T203 : ex_ra3;
  assign T203 = io_inst[5'h18:5'h14];
  assign T204 = T205 & fp_decoder_io_sigs_swap23;
  assign T205 = io_valid & fp_decoder_io_sigs_ren2;
  assign T206 = io_inst[5'h1f:5'h1b];
  assign T207 = io_valid & fp_decoder_io_sigs_ren3;
  assign req_in2 = T208;
  assign T208 = ex_reg_valid ? ex_rs2 : cp_rs2;
  assign cp_rs2 = io_cp_req_bits_swap23 ? io_cp_req_bits_in3 : io_cp_req_bits_in2;
  assign ex_rs2 = regfile[ex_ra2];
  assign T209 = T215 ? T214 : T210;
  assign T210 = T212 ? T211 : ex_ra2;
  assign T211 = io_inst[5'h13:4'hf];
  assign T212 = T213 & fp_decoder_io_sigs_swap12;
  assign T213 = io_valid & fp_decoder_io_sigs_ren1;
  assign T214 = io_inst[5'h18:5'h14];
  assign T215 = T205 & T216;
  assign T216 = T218 & T217;
  assign T217 = fp_decoder_io_sigs_swap23 ^ 1'h1;
  assign T218 = fp_decoder_io_sigs_swap12 ^ 1'h1;
  assign req_in1 = T219;
  assign T219 = ex_reg_valid ? ex_rs1 : io_cp_req_bits_in1;
  assign ex_rs1 = regfile[ex_ra1];
  assign T220 = T226 ? T225 : T221;
  assign T221 = T223 ? T222 : ex_ra1;
  assign T222 = io_inst[5'h13:4'hf];
  assign T223 = T213 & T224;
  assign T224 = fp_decoder_io_sigs_swap12 ^ 1'h1;
  assign T225 = io_inst[5'h18:5'h14];
  assign T226 = T205 & fp_decoder_io_sigs_swap12;
  assign req_typ = T227;
  assign T227 = ex_reg_valid ? T228 : io_cp_req_bits_typ;
  assign T228 = ex_reg_inst[5'h15:5'h14];
  assign req_rm = T229;
  assign T229 = ex_reg_valid ? ex_rm : io_cp_req_bits_rm;
  assign ex_rm = T231 ? io_fcsr_rm : T230;
  assign T230 = ex_reg_inst[4'he:4'hc];
  assign T231 = T232 == 3'h7;
  assign T232 = ex_reg_inst[4'he:4'hc];
  assign req_wflags = T233;
  assign T233 = ex_reg_valid ? R234 : cp_ctrl_wflags;
  assign cp_ctrl_wflags = io_cp_req_bits_wflags;
  assign T235 = io_valid ? fp_decoder_io_sigs_wflags : R234;
  assign req_round = T236;
  assign T236 = ex_reg_valid ? R237 : cp_ctrl_round;
  assign cp_ctrl_round = io_cp_req_bits_round;
  assign T238 = io_valid ? fp_decoder_io_sigs_round : R237;
  assign req_sqrt = T8;
  assign req_div = T18;
  assign req_fma = T45;
  assign req_fastpipe = T57;
  assign req_toint = T239;
  assign T239 = ex_reg_valid ? R240 : cp_ctrl_toint;
  assign cp_ctrl_toint = io_cp_req_bits_toint;
  assign T241 = io_valid ? fp_decoder_io_sigs_toint : R240;
  assign req_fromint = T53;
  assign req_single = T41;
  assign req_swap23 = T242;
  assign T242 = ex_reg_valid ? R243 : cp_ctrl_swap23;
  assign cp_ctrl_swap23 = io_cp_req_bits_swap23;
  assign T244 = io_valid ? fp_decoder_io_sigs_swap23 : R243;
  assign req_swap12 = T245;
  assign T245 = ex_reg_valid ? R246 : cp_ctrl_swap12;
  assign cp_ctrl_swap12 = io_cp_req_bits_swap12;
  assign T247 = io_valid ? fp_decoder_io_sigs_swap12 : R246;
  assign req_ren3 = T248;
  assign T248 = ex_reg_valid ? R249 : cp_ctrl_ren3;
  assign cp_ctrl_ren3 = io_cp_req_bits_ren3;
  assign T250 = io_valid ? fp_decoder_io_sigs_ren3 : R249;
  assign req_ren2 = T251;
  assign T251 = ex_reg_valid ? R252 : cp_ctrl_ren2;
  assign cp_ctrl_ren2 = io_cp_req_bits_ren2;
  assign T253 = io_valid ? fp_decoder_io_sigs_ren2 : R252;
  assign req_ren1 = T254;
  assign T254 = ex_reg_valid ? R255 : cp_ctrl_ren1;
  assign cp_ctrl_ren1 = io_cp_req_bits_ren1;
  assign T256 = io_valid ? fp_decoder_io_sigs_ren1 : R255;
  assign req_wen = T257;
  assign T257 = ex_reg_valid ? R258 : cp_ctrl_wen;
  assign cp_ctrl_wen = io_cp_req_bits_wen;
  assign T259 = io_valid ? fp_decoder_io_sigs_wen : R258;
  assign req_ldst = T260;
  assign T260 = ex_reg_valid ? R261 : cp_ctrl_ldst;
  assign cp_ctrl_ldst = io_cp_req_bits_ldst;
  assign T262 = io_valid ? fp_decoder_io_sigs_ldst : R261;
  assign req_cmd = T263;
  assign T263 = ex_reg_valid ? R264 : cp_ctrl_cmd;
  assign cp_ctrl_cmd = io_cp_req_bits_cmd;
  assign T265 = io_valid ? fp_decoder_io_sigs_cmd : R264;
  assign T266 = req_valid & T57;
  assign T267 = ex_reg_valid ? T556 : io_cp_req_bits_in1;
  assign T556 = {1'h0, io_fromint_data};
  assign T268 = req_valid & T53;
  assign T269 = req_valid & T270;
  assign T270 = T273 | T271;
  assign T271 = 5'h5 == T272;
  assign T272 = T263 & 5'hd;
  assign T273 = T274 | T8;
  assign T274 = T239 | T18;
  assign T275 = T277 & T276;
  assign T276 = T41 ^ 1'h1;
  assign T277 = req_valid & T45;
  assign T278 = T279 & T41;
  assign T279 = req_valid & T45;
  assign io_cp_resp_bits_data = T280;
  assign T280 = T285 ? wdata : T557;
  assign T557 = {1'h0, T281};
  assign T281 = T282 ? fpiu_io_out_bits_toint : 64'h0;
  assign T282 = T284 & mem_ctrl_toint;
  assign T283 = req_valid ? T239 : mem_ctrl_toint;
  assign T284 = fpiu_io_out_valid & mem_cp_valid;
  assign T285 = wcp & T286;
  assign T286 = wen[1'h0];
  assign io_cp_resp_valid = T287;
  assign T287 = T285 ? 1'h1 : T282;
  assign io_cp_req_ready = T288;
  assign T288 = ex_reg_valid ^ 1'h1;
  assign io_sboard_clra = waddr;
  assign io_sboard_clr = T289;
  assign T289 = T290 & divSqrt_wen;
  assign T290 = wb_cp_valid ^ 1'h1;
  assign T558 = reset ? 1'h0 : mem_cp_valid;
  assign io_sboard_set = T291;
  assign T291 = T294 & R292;
  assign T293 = mem_ctrl_div | mem_ctrl_sqrt;
  assign T294 = wb_reg_valid & T295;
  assign T295 = wb_cp_valid ^ 1'h1;
  assign T559 = reset ? 1'h0 : T296;
  assign T296 = mem_reg_valid & T297;
  assign T297 = T298 | mem_cp_valid;
  assign T298 = killm ^ 1'h1;
  assign io_dec_wflags = fp_decoder_io_sigs_wflags;
  assign io_dec_round = fp_decoder_io_sigs_round;
  assign io_dec_sqrt = fp_decoder_io_sigs_sqrt;
  assign io_dec_div = fp_decoder_io_sigs_div;
  assign io_dec_fma = fp_decoder_io_sigs_fma;
  assign io_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_dec_toint = fp_decoder_io_sigs_toint;
  assign io_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_dec_single = fp_decoder_io_sigs_single;
  assign io_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_dec_swap12 = fp_decoder_io_sigs_swap12;
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_dec_wen = fp_decoder_io_sigs_wen;
  assign io_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_illegal_rm = T299;
  assign T299 = T300 & T236;
  assign T300 = ex_rm[2'h2];
  assign io_nack_mem = T301;
  assign T301 = T302 | divSqrt_in_flight;
  assign T302 = units_busy | write_port_busy;
  assign units_busy = T306 & T303;
  assign T303 = T305 | T304;
  assign T304 = wen != 2'h0;
  assign T305 = divSqrt_inReady ^ 1'h1;
  assign T306 = mem_reg_valid & T307;
  assign T307 = mem_ctrl_div | mem_ctrl_sqrt;
  assign io_fcsr_rdy = T308;
  assign T308 = T309 ^ 1'h1;
  assign T309 = T310 | divSqrt_in_flight;
  assign T310 = T312 | T311;
  assign T311 = wen != 2'h0;
  assign T312 = T315 | T313;
  assign T313 = wb_reg_valid & wb_ctrl_toint;
  assign T314 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign T315 = T318 | T316;
  assign T316 = mem_reg_valid & mem_ctrl_wflags;
  assign T317 = req_valid ? T233 : mem_ctrl_wflags;
  assign T318 = ex_reg_valid & T233;
  assign io_toint_data = fpiu_io_out_bits_toint;
  assign io_store_data = fpiu_io_out_bits_store;
  assign io_fcsr_flags_bits = T319;
  assign T319 = T328 | T320;
  assign T320 = T327 ? wexc : 5'h0;
  assign wexc = T326 ? T324 : T321;
  assign T321 = T322 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign T322 = T323[1'h0];
  assign T323 = T560;
  assign T560 = wsrc[1'h1:1'h0];
  assign T324 = T325 ? dfma_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T325 = T323[1'h0];
  assign T326 = T323[1'h1];
  assign T327 = wen[1'h0];
  assign T328 = T334 | T329;
  assign T329 = divSqrt_wen ? divSqrt_flags : 5'h0;
  assign divSqrt_flags = T330;
  assign T330 = R332 | T331;
  assign T331 = R120 ? RecFNToRecFN_io_exceptionFlags : 5'h0;
  assign T333 = T6 ? DivSqrtRecF64_io_exceptionFlags : R332;
  assign T334 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T335 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign io_fcsr_flags_valid = T336;
  assign T336 = T338 | T337;
  assign T337 = wen[1'h0];
  assign T338 = wb_toint_valid | divSqrt_wen;
  FPUDecoder fp_decoder(
       .io_inst( io_inst ),
       .io_sigs_cmd( fp_decoder_io_sigs_cmd ),
       .io_sigs_ldst( fp_decoder_io_sigs_ldst ),
       .io_sigs_wen( fp_decoder_io_sigs_wen ),
       .io_sigs_ren1( fp_decoder_io_sigs_ren1 ),
       .io_sigs_ren2( fp_decoder_io_sigs_ren2 ),
       .io_sigs_ren3( fp_decoder_io_sigs_ren3 ),
       .io_sigs_swap12( fp_decoder_io_sigs_swap12 ),
       .io_sigs_swap23( fp_decoder_io_sigs_swap23 ),
       .io_sigs_single( fp_decoder_io_sigs_single ),
       .io_sigs_fromint( fp_decoder_io_sigs_fromint ),
       .io_sigs_toint( fp_decoder_io_sigs_toint ),
       .io_sigs_fastpipe( fp_decoder_io_sigs_fastpipe ),
       .io_sigs_fma( fp_decoder_io_sigs_fma ),
       .io_sigs_div( fp_decoder_io_sigs_div ),
       .io_sigs_sqrt( fp_decoder_io_sigs_sqrt ),
       .io_sigs_round( fp_decoder_io_sigs_round ),
       .io_sigs_wflags( fp_decoder_io_sigs_wflags )
  );
  FPUFMAPipe_0 sfma(.clk(clk), .reset(reset),
       .io_in_valid( T278 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap12( req_swap12 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_div( req_div ),
       .io_in_bits_sqrt( req_sqrt ),
       .io_in_bits_round( req_round ),
       .io_in_bits_wflags( req_wflags ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( sfma_io_out_bits_data ),
       .io_out_bits_exc( sfma_io_out_bits_exc )
  );
  FPUFMAPipe_1 dfma(.clk(clk), .reset(reset),
       .io_in_valid( T275 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap12( req_swap12 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_div( req_div ),
       .io_in_bits_sqrt( req_sqrt ),
       .io_in_bits_round( req_round ),
       .io_in_bits_wflags( req_wflags ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( dfma_io_out_bits_data ),
       .io_out_bits_exc( dfma_io_out_bits_exc )
  );
  FPToInt fpiu(.clk(clk),
       .io_in_valid( T269 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap12( req_swap12 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_div( req_div ),
       .io_in_bits_sqrt( req_sqrt ),
       .io_in_bits_round( req_round ),
       .io_in_bits_wflags( req_wflags ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_as_double_cmd(  )
       //.io_as_double_ldst(  )
       //.io_as_double_wen(  )
       //.io_as_double_ren1(  )
       //.io_as_double_ren2(  )
       //.io_as_double_ren3(  )
       //.io_as_double_swap12(  )
       //.io_as_double_swap23(  )
       //.io_as_double_single(  )
       //.io_as_double_fromint(  )
       //.io_as_double_toint(  )
       //.io_as_double_fastpipe(  )
       //.io_as_double_fma(  )
       //.io_as_double_div(  )
       //.io_as_double_sqrt(  )
       //.io_as_double_round(  )
       //.io_as_double_wflags(  )
       .io_as_double_rm( fpiu_io_as_double_rm ),
       //.io_as_double_typ(  )
       .io_as_double_in1( fpiu_io_as_double_in1 ),
       .io_as_double_in2( fpiu_io_as_double_in2 ),
       //.io_as_double_in3(  )
       .io_out_valid( fpiu_io_out_valid ),
       .io_out_bits_lt( fpiu_io_out_bits_lt ),
       .io_out_bits_store( fpiu_io_out_bits_store ),
       .io_out_bits_toint( fpiu_io_out_bits_toint ),
       .io_out_bits_exc( fpiu_io_out_bits_exc )
  );
  IntToFP ifpu(.clk(clk), .reset(reset),
       .io_in_valid( T268 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap12( req_swap12 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_div( req_div ),
       .io_in_bits_sqrt( req_sqrt ),
       .io_in_bits_round( req_round ),
       .io_in_bits_wflags( req_wflags ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( T267 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( ifpu_io_out_bits_data ),
       .io_out_bits_exc( ifpu_io_out_bits_exc )
  );
  FPToFP fpmu(.clk(clk), .reset(reset),
       .io_in_valid( T266 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap12( req_swap12 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_div( req_div ),
       .io_in_bits_sqrt( req_sqrt ),
       .io_in_bits_round( req_round ),
       .io_in_bits_wflags( req_wflags ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( fpmu_io_out_bits_data ),
       .io_out_bits_exc( fpmu_io_out_bits_exc ),
       .io_lt( fpiu_io_out_bits_lt )
  );
  DivSqrtRecF64 DivSqrtRecF64(.clk(clk), .reset(reset),
       .io_inReady_div( DivSqrtRecF64_io_inReady_div ),
       .io_inReady_sqrt( DivSqrtRecF64_io_inReady_sqrt ),
       .io_inValid( T11 ),
       .io_sqrtOp( mem_ctrl_sqrt ),
       .io_a( fpiu_io_as_double_in1 ),
       .io_b( fpiu_io_as_double_in2 ),
       .io_roundingMode( T339 ),
       .io_outValid_div( DivSqrtRecF64_io_outValid_div ),
       .io_outValid_sqrt( DivSqrtRecF64_io_outValid_sqrt ),
       .io_out( DivSqrtRecF64_io_out ),
       .io_exceptionFlags( DivSqrtRecF64_io_exceptionFlags )
  );
  RecFNToRecFN_1 RecFNToRecFN(
       .io_in( R4 ),
       .io_roundingMode( R0 ),
       .io_out( RecFNToRecFN_io_out ),
       .io_exceptionFlags( RecFNToRecFN_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(T2) begin
      R0 <= T339;
    end
    if(T6) begin
      R4 <= DivSqrtRecF64_io_out;
    end
    if(req_valid) begin
      mem_ctrl_sqrt <= T8;
    end
    if(io_valid) begin
      R9 <= fp_decoder_io_sigs_sqrt;
    end
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if(reset) begin
      divSqrt_in_flight <= 1'h0;
    end else if(T6) begin
      divSqrt_in_flight <= 1'h0;
    end else if(T2) begin
      divSqrt_in_flight <= 1'h1;
    end
    if(req_valid) begin
      mem_ctrl_div <= T18;
    end
    if(io_valid) begin
      R19 <= fp_decoder_io_sigs_div;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T21;
    end
    if (T125)
      regfile[waddr] <= wdata;
    if(T112) begin
      winfo_0 <= mem_winfo;
    end else if(T98) begin
      winfo_0 <= winfo_1;
    end
    if(T34) begin
      winfo_1 <= mem_winfo;
    end
    if(req_valid) begin
      mem_ctrl_single <= T41;
    end
    if(io_valid) begin
      R42 <= fp_decoder_io_sigs_single;
    end
    if(req_valid) begin
      mem_ctrl_fma <= T45;
    end
    if(io_valid) begin
      R46 <= fp_decoder_io_sigs_fma;
    end
    if(req_valid) begin
      mem_ctrl_fromint <= T53;
    end
    if(io_valid) begin
      R54 <= fp_decoder_io_sigs_fromint;
    end
    if(req_valid) begin
      mem_ctrl_fastpipe <= T57;
    end
    if(io_valid) begin
      R58 <= fp_decoder_io_sigs_fastpipe;
    end
    if(req_valid) begin
      write_port_busy <= T62;
    end
    if(reset) begin
      wen <= 2'h0;
    end else if(T79) begin
      wen <= T77;
    end else begin
      wen <= T350;
    end
    if(reset) begin
      mem_cp_valid <= 1'h0;
    end else begin
      mem_cp_valid <= ex_cp_valid;
    end
    if(ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(io_valid) begin
      ex_reg_inst <= io_inst;
    end
    if(T2) begin
      R120 <= mem_ctrl_single;
    end
    if(T6) begin
      divSqrt_wen <= T123;
    end else begin
      divSqrt_wen <= 1'h0;
    end
    if(T2) begin
      divSqrt_killed <= killm;
    end
    if(T2) begin
      divSqrt_waddr <= T132;
    end
    if (load_wb)
      regfile[load_wb_tag] <= load_wb_data_recoded;
    if(io_dmem_resp_val) begin
      load_wb_data <= io_dmem_resp_data;
    end
    if(io_dmem_resp_val) begin
      load_wb_single <= T197;
    end
    load_wb <= io_dmem_resp_val;
    if(io_dmem_resp_val) begin
      load_wb_tag <= io_dmem_resp_tag;
    end
    if(T207) begin
      ex_ra3 <= T206;
    end else if(T204) begin
      ex_ra3 <= T203;
    end
    if(T215) begin
      ex_ra2 <= T214;
    end else if(T212) begin
      ex_ra2 <= T211;
    end
    if(T226) begin
      ex_ra1 <= T225;
    end else if(T223) begin
      ex_ra1 <= T222;
    end
    if(io_valid) begin
      R234 <= fp_decoder_io_sigs_wflags;
    end
    if(io_valid) begin
      R237 <= fp_decoder_io_sigs_round;
    end
    if(io_valid) begin
      R240 <= fp_decoder_io_sigs_toint;
    end
    if(io_valid) begin
      R243 <= fp_decoder_io_sigs_swap23;
    end
    if(io_valid) begin
      R246 <= fp_decoder_io_sigs_swap12;
    end
    if(io_valid) begin
      R249 <= fp_decoder_io_sigs_ren3;
    end
    if(io_valid) begin
      R252 <= fp_decoder_io_sigs_ren2;
    end
    if(io_valid) begin
      R255 <= fp_decoder_io_sigs_ren1;
    end
    if(io_valid) begin
      R258 <= fp_decoder_io_sigs_wen;
    end
    if(io_valid) begin
      R261 <= fp_decoder_io_sigs_ldst;
    end
    if(io_valid) begin
      R264 <= fp_decoder_io_sigs_cmd;
    end
    if(req_valid) begin
      mem_ctrl_toint <= T239;
    end
    if(reset) begin
      wb_cp_valid <= 1'h0;
    end else begin
      wb_cp_valid <= mem_cp_valid;
    end
    R292 <= T293;
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T296;
    end
    if(mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if(req_valid) begin
      mem_ctrl_wflags <= T233;
    end
    if(T6) begin
      R332 <= DivSqrtRecF64_io_exceptionFlags;
    end
    if(mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [5:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [5:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[5:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T54;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T55;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  locked;
  wire T56;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  reg [1:0] R20;
  wire[1:0] T57;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[127:0] T24;
  wire T25;
  wire[16:0] T26;
  wire[2:0] T27;
  wire T28;
  wire[1:0] T29;
  wire[5:0] T30;
  wire[25:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T54 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T55 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T14 & T12;
  assign T12 = io_out_bits_is_builtin_type & T13;
  assign T13 = 3'h3 == io_out_bits_a_type;
  assign T14 = io_out_valid & io_out_ready;
  assign T56 = reset ? 1'h0 : T15;
  assign T15 = T22 ? 1'h0 : T16;
  assign T16 = T11 ? T17 : locked;
  assign T17 = T18 ^ 1'h1;
  assign T18 = T19 == 2'h0;
  assign T19 = R20 + 2'h1;
  assign T57 = reset ? 2'h0 : T21;
  assign T21 = T11 ? T19 : R20;
  assign T22 = T14 & T23;
  assign T23 = T12 ^ 1'h1;
  assign io_out_bits_data = T24;
  assign T24 = T25 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T25 = chosen;
  assign io_out_bits_union = T26;
  assign T26 = T25 ? io_in_1_bits_union : io_in_0_bits_union;
  assign io_out_bits_a_type = T27;
  assign T27 = T25 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_is_builtin_type = T28;
  assign T28 = T25 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_addr_beat = T29;
  assign T29 = T25 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T30;
  assign T30 = T25 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T31;
  assign T31 = T25 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T32;
  assign T32 = T25 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T33;
  assign T33 = T34 & io_out_ready;
  assign T34 = locked ? T43 : T35;
  assign T35 = T42 | T36;
  assign T36 = T37 ^ 1'h1;
  assign T37 = T40 | T38;
  assign T38 = io_in_1_valid & T39;
  assign T39 = last_grant < 1'h1;
  assign T40 = io_in_0_valid & T41;
  assign T41 = last_grant < 1'h0;
  assign T42 = last_grant < 1'h0;
  assign T43 = lockIdx == 1'h0;
  assign io_in_1_ready = T44;
  assign T44 = T45 & io_out_ready;
  assign T45 = locked ? T53 : T46;
  assign T46 = T50 | T47;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_0_valid;
  assign T49 = T40 | T38;
  assign T50 = T52 & T51;
  assign T51 = last_grant < 1'h1;
  assign T52 = T40 ^ 1'h1;
  assign T53 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T22) begin
      locked <= 1'h0;
    end else if(T11) begin
      locked <= T17;
    end
    if(reset) begin
      R20 <= 2'h0;
    end else if(T11) begin
      R20 <= T19;
    end
  end
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [5:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_voluntary,
    input [2:0] io_in_1_bits_r_type,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [5:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_voluntary,
    input [2:0] io_in_0_bits_r_type,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[5:0] io_out_bits_client_xact_id,
    output io_out_bits_voluntary,
    output[2:0] io_out_bits_r_type,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T56;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T57;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  locked;
  wire T58;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  reg [1:0] R23;
  wire[1:0] T59;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[127:0] T27;
  wire T28;
  wire[2:0] T29;
  wire T30;
  wire[5:0] T31;
  wire[25:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R23 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T56 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T57 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T17 & T12;
  assign T12 = T14 | T13;
  assign T13 = 3'h2 == io_out_bits_r_type;
  assign T14 = T16 | T15;
  assign T15 = 3'h1 == io_out_bits_r_type;
  assign T16 = 3'h0 == io_out_bits_r_type;
  assign T17 = io_out_valid & io_out_ready;
  assign T58 = reset ? 1'h0 : T18;
  assign T18 = T25 ? 1'h0 : T19;
  assign T19 = T11 ? T20 : locked;
  assign T20 = T21 ^ 1'h1;
  assign T21 = T22 == 2'h0;
  assign T22 = R23 + 2'h1;
  assign T59 = reset ? 2'h0 : T24;
  assign T24 = T11 ? T22 : R23;
  assign T25 = T17 & T26;
  assign T26 = T12 ^ 1'h1;
  assign io_out_bits_data = T27;
  assign T27 = T28 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T28 = chosen;
  assign io_out_bits_r_type = T29;
  assign T29 = T28 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_voluntary = T30;
  assign T30 = T28 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_client_xact_id = T31;
  assign T31 = T28 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T32;
  assign T32 = T28 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T33;
  assign T33 = T28 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T34;
  assign T34 = T28 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T35;
  assign T35 = T36 & io_out_ready;
  assign T36 = locked ? T45 : T37;
  assign T37 = T44 | T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T42 | T40;
  assign T40 = io_in_1_valid & T41;
  assign T41 = last_grant < 1'h1;
  assign T42 = io_in_0_valid & T43;
  assign T43 = last_grant < 1'h0;
  assign T44 = last_grant < 1'h0;
  assign T45 = lockIdx == 1'h0;
  assign io_in_1_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = locked ? T55 : T48;
  assign T48 = T52 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_0_valid;
  assign T51 = T42 | T40;
  assign T52 = T54 & T53;
  assign T53 = last_grant < 1'h1;
  assign T54 = T42 ^ 1'h1;
  assign T55 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T25) begin
      locked <= 1'h0;
    end else if(T11) begin
      locked <= T20;
    end
    if(reset) begin
      R23 <= 2'h0;
    end else if(T11) begin
      R23 <= T22;
    end
  end
endmodule

module ClientTileLinkIOArbiter(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [25:0] io_in_1_acquire_bits_addr_block,
    input [5:0] io_in_1_acquire_bits_client_xact_id,
    input [1:0] io_in_1_acquire_bits_addr_beat,
    input  io_in_1_acquire_bits_is_builtin_type,
    input [2:0] io_in_1_acquire_bits_a_type,
    input [16:0] io_in_1_acquire_bits_union,
    input [127:0] io_in_1_acquire_bits_data,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_addr_beat,
    output[5:0] io_in_1_grant_bits_client_xact_id,
    output[3:0] io_in_1_grant_bits_manager_xact_id,
    output io_in_1_grant_bits_is_builtin_type,
    output[3:0] io_in_1_grant_bits_g_type,
    output[127:0] io_in_1_grant_bits_data,
    input  io_in_1_probe_ready,
    output io_in_1_probe_valid,
    output[25:0] io_in_1_probe_bits_addr_block,
    output[1:0] io_in_1_probe_bits_p_type,
    output io_in_1_release_ready,
    input  io_in_1_release_valid,
    input [1:0] io_in_1_release_bits_addr_beat,
    input [25:0] io_in_1_release_bits_addr_block,
    input [5:0] io_in_1_release_bits_client_xact_id,
    input  io_in_1_release_bits_voluntary,
    input [2:0] io_in_1_release_bits_r_type,
    input [127:0] io_in_1_release_bits_data,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [25:0] io_in_0_acquire_bits_addr_block,
    input [5:0] io_in_0_acquire_bits_client_xact_id,
    input [1:0] io_in_0_acquire_bits_addr_beat,
    input  io_in_0_acquire_bits_is_builtin_type,
    input [2:0] io_in_0_acquire_bits_a_type,
    input [16:0] io_in_0_acquire_bits_union,
    input [127:0] io_in_0_acquire_bits_data,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_addr_beat,
    output[5:0] io_in_0_grant_bits_client_xact_id,
    output[3:0] io_in_0_grant_bits_manager_xact_id,
    output io_in_0_grant_bits_is_builtin_type,
    output[3:0] io_in_0_grant_bits_g_type,
    output[127:0] io_in_0_grant_bits_data,
    input  io_in_0_probe_ready,
    output io_in_0_probe_valid,
    output[25:0] io_in_0_probe_bits_addr_block,
    output[1:0] io_in_0_probe_bits_p_type,
    output io_in_0_release_ready,
    input  io_in_0_release_valid,
    input [1:0] io_in_0_release_bits_addr_beat,
    input [25:0] io_in_0_release_bits_addr_block,
    input [5:0] io_in_0_release_bits_client_xact_id,
    input  io_in_0_release_bits_voluntary,
    input [2:0] io_in_0_release_bits_r_type,
    input [127:0] io_in_0_release_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[5:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [5:0] io_out_grant_bits_client_xact_id,
    input [3:0] io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid,
    output[1:0] io_out_release_bits_addr_beat,
    output[25:0] io_out_release_bits_addr_block,
    output[5:0] io_out_release_bits_client_xact_id,
    output io_out_release_bits_voluntary,
    output[2:0] io_out_release_bits_r_type,
    output[127:0] io_out_release_bits_data
);

  wire[5:0] T17;
  wire[6:0] T0;
  wire[5:0] T18;
  wire[6:0] T1;
  wire[5:0] T19;
  wire[6:0] T2;
  wire[5:0] T20;
  wire[6:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[5:0] T21;
  wire[4:0] T13;
  wire T14;
  wire[5:0] T22;
  wire[4:0] T15;
  wire T16;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[25:0] LockingRRArbiter_io_out_bits_addr_block;
  wire[5:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_addr_beat;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_union;
  wire[127:0] LockingRRArbiter_io_out_bits_data;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_addr_beat;
  wire[25:0] LockingRRArbiter_1_io_out_bits_addr_block;
  wire[5:0] LockingRRArbiter_1_io_out_bits_client_xact_id;
  wire LockingRRArbiter_1_io_out_bits_voluntary;
  wire[2:0] LockingRRArbiter_1_io_out_bits_r_type;
  wire[127:0] LockingRRArbiter_1_io_out_bits_data;


  assign T17 = T0[3'h5:1'h0];
  assign T0 = {io_in_0_release_bits_client_xact_id, 1'h0};
  assign T18 = T1[3'h5:1'h0];
  assign T1 = {io_in_1_release_bits_client_xact_id, 1'h1};
  assign T19 = T2[3'h5:1'h0];
  assign T2 = {io_in_0_acquire_bits_client_xact_id, 1'h0};
  assign T20 = T3[3'h5:1'h0];
  assign T3 = {io_in_1_acquire_bits_client_xact_id, 1'h1};
  assign io_out_release_bits_data = LockingRRArbiter_1_io_out_bits_data;
  assign io_out_release_bits_r_type = LockingRRArbiter_1_io_out_bits_r_type;
  assign io_out_release_bits_voluntary = LockingRRArbiter_1_io_out_bits_voluntary;
  assign io_out_release_bits_client_xact_id = LockingRRArbiter_1_io_out_bits_client_xact_id;
  assign io_out_release_bits_addr_block = LockingRRArbiter_1_io_out_bits_addr_block;
  assign io_out_release_bits_addr_beat = LockingRRArbiter_1_io_out_bits_addr_beat;
  assign io_out_release_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_probe_ready = T4;
  assign T4 = io_in_0_probe_ready & io_in_1_probe_ready;
  assign io_out_grant_ready = T5;
  assign T5 = T10 ? io_in_1_grant_ready : T6;
  assign T6 = T7 ? io_in_0_grant_ready : 1'h0;
  assign T7 = T8 == 1'h0;
  assign T8 = T9;
  assign T9 = io_out_grant_bits_client_xact_id[1'h0];
  assign T10 = T11 == 1'h1;
  assign T11 = T12;
  assign T12 = io_out_grant_bits_client_xact_id[1'h0];
  assign io_out_acquire_bits_data = LockingRRArbiter_io_out_bits_data;
  assign io_out_acquire_bits_union = LockingRRArbiter_io_out_bits_union;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_io_out_bits_addr_block;
  assign io_out_acquire_valid = LockingRRArbiter_io_out_valid;
  assign io_in_0_release_ready = LockingRRArbiter_1_io_in_0_ready;
  assign io_in_0_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_0_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_0_probe_valid = io_out_probe_valid;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_client_xact_id = T21;
  assign T21 = {1'h0, T13};
  assign T13 = io_out_grant_bits_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_valid = T14;
  assign T14 = T7 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_io_in_0_ready;
  assign io_in_1_release_ready = LockingRRArbiter_1_io_in_1_ready;
  assign io_in_1_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_1_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_1_probe_valid = io_out_probe_valid;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_client_xact_id = T22;
  assign T22 = {1'h0, T15};
  assign T15 = io_out_grant_bits_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_valid = T16;
  assign T16 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_io_in_1_ready;
  LockingRRArbiter_0 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_addr_block( io_in_1_acquire_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T20 ),
       .io_in_1_bits_addr_beat( io_in_1_acquire_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( io_in_1_acquire_bits_is_builtin_type ),
       .io_in_1_bits_a_type( io_in_1_acquire_bits_a_type ),
       .io_in_1_bits_union( io_in_1_acquire_bits_union ),
       .io_in_1_bits_data( io_in_1_acquire_bits_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_addr_block( io_in_0_acquire_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T19 ),
       .io_in_0_bits_addr_beat( io_in_0_acquire_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( io_in_0_acquire_bits_is_builtin_type ),
       .io_in_0_bits_a_type( io_in_0_acquire_bits_a_type ),
       .io_in_0_bits_union( io_in_0_acquire_bits_union ),
       .io_in_0_bits_data( io_in_0_acquire_bits_data ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( LockingRRArbiter_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( LockingRRArbiter_io_out_bits_a_type ),
       .io_out_bits_union( LockingRRArbiter_io_out_bits_union ),
       .io_out_bits_data( LockingRRArbiter_io_out_bits_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_release_valid ),
       .io_in_1_bits_addr_beat( io_in_1_release_bits_addr_beat ),
       .io_in_1_bits_addr_block( io_in_1_release_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T18 ),
       .io_in_1_bits_voluntary( io_in_1_release_bits_voluntary ),
       .io_in_1_bits_r_type( io_in_1_release_bits_r_type ),
       .io_in_1_bits_data( io_in_1_release_bits_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_release_valid ),
       .io_in_0_bits_addr_beat( io_in_0_release_bits_addr_beat ),
       .io_in_0_bits_addr_block( io_in_0_release_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T17 ),
       .io_in_0_bits_voluntary( io_in_0_release_bits_voluntary ),
       .io_in_0_bits_r_type( io_in_0_release_bits_r_type ),
       .io_in_0_bits_data( io_in_0_release_bits_data ),
       .io_out_ready( io_out_release_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_addr_beat( LockingRRArbiter_1_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( LockingRRArbiter_1_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_1_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( LockingRRArbiter_1_io_out_bits_voluntary ),
       .io_out_bits_r_type( LockingRRArbiter_1_io_out_bits_r_type ),
       .io_out_bits_data( LockingRRArbiter_1_io_out_bits_data )
       //.io_chosen(  )
  );
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [4:0] io_in_0_bits_rd,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[4:0] io_out_bits_rd,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_rd = io_in_0_bits_rd;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [6:0] io_enq_bits_inst_funct,
    input [4:0] io_enq_bits_inst_rs2,
    input [4:0] io_enq_bits_inst_rs1,
    input  io_enq_bits_inst_xd,
    input  io_enq_bits_inst_xs1,
    input  io_enq_bits_inst_xs2,
    input [4:0] io_enq_bits_inst_rd,
    input [6:0] io_enq_bits_inst_opcode,
    input [63:0] io_enq_bits_rs1,
    input [63:0] io_enq_bits_rs2,
    input  io_deq_ready,
    output io_deq_valid,
    output[6:0] io_deq_bits_inst_funct,
    output[4:0] io_deq_bits_inst_rs2,
    output[4:0] io_deq_bits_inst_rs1,
    output io_deq_bits_inst_xd,
    output io_deq_bits_inst_xs1,
    output io_deq_bits_inst_xs2,
    output[4:0] io_deq_bits_inst_rd,
    output[6:0] io_deq_bits_inst_opcode,
    output[63:0] io_deq_bits_rs1,
    output[63:0] io_deq_bits_rs2,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T35;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T36;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T37;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[159:0] T11;
  reg [159:0] ram [1:0];
  wire[159:0] T12;
  wire[159:0] T13;
  wire[159:0] T14;
  wire[140:0] T15;
  wire[134:0] T16;
  wire[127:0] T17;
  wire[5:0] T18;
  wire[18:0] T19;
  wire[6:0] T20;
  wire[1:0] T21;
  wire[11:0] T22;
  wire[63:0] T23;
  wire[6:0] T24;
  wire[4:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[4:0] T29;
  wire[4:0] T30;
  wire[6:0] T31;
  wire T32;
  wire empty;
  wire T33;
  wire T34;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T35 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T36 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T37 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rs2 = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T19, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_inst_opcode, T17};
  assign T17 = {io_enq_bits_rs1, io_enq_bits_rs2};
  assign T18 = {io_enq_bits_inst_xs2, io_enq_bits_inst_rd};
  assign T19 = {T22, T20};
  assign T20 = {io_enq_bits_inst_rs1, T21};
  assign T21 = {io_enq_bits_inst_xd, io_enq_bits_inst_xs1};
  assign T22 = {io_enq_bits_inst_funct, io_enq_bits_inst_rs2};
  assign io_deq_bits_rs1 = T23;
  assign T23 = T11[7'h7f:7'h40];
  assign io_deq_bits_inst_opcode = T24;
  assign T24 = T11[8'h86:8'h80];
  assign io_deq_bits_inst_rd = T25;
  assign T25 = T11[8'h8b:8'h87];
  assign io_deq_bits_inst_xs2 = T26;
  assign T26 = T11[8'h8c];
  assign io_deq_bits_inst_xs1 = T27;
  assign T27 = T11[8'h8d];
  assign io_deq_bits_inst_xd = T28;
  assign T28 = T11[8'h8e];
  assign io_deq_bits_inst_rs1 = T29;
  assign T29 = T11[8'h93:8'h8f];
  assign io_deq_bits_inst_rs2 = T30;
  assign T30 = T11[8'h98:8'h94];
  assign io_deq_bits_inst_funct = T31;
  assign T31 = T11[8'h9f:8'h99];
  assign io_deq_valid = T32;
  assign T32 = empty ^ 1'h1;
  assign empty = ptr_match & T33;
  assign T33 = maybe_full ^ 1'h1;
  assign io_enq_ready = T34;
  assign T34 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module RoccCommandRouter(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [6:0] io_in_bits_inst_funct,
    input [4:0] io_in_bits_inst_rs2,
    input [4:0] io_in_bits_inst_rs1,
    input  io_in_bits_inst_xd,
    input  io_in_bits_inst_xs1,
    input  io_in_bits_inst_xs2,
    input [4:0] io_in_bits_inst_rd,
    input [6:0] io_in_bits_inst_opcode,
    input [63:0] io_in_bits_rs1,
    input [63:0] io_in_bits_rs2,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[6:0] io_out_0_bits_inst_funct,
    output[4:0] io_out_0_bits_inst_rs2,
    output[4:0] io_out_0_bits_inst_rs1,
    output io_out_0_bits_inst_xd,
    output io_out_0_bits_inst_xs1,
    output io_out_0_bits_inst_xs2,
    output[4:0] io_out_0_bits_inst_rd,
    output[6:0] io_out_0_bits_inst_opcode,
    output[63:0] io_out_0_bits_rs1,
    output[63:0] io_out_0_bits_rs2,
    output io_busy
);

  reg  T0;
  wire T1;
  wire T2;
  wire cmdReadys_0;
  wire T3;
  wire T4;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[6:0] Queue_io_deq_bits_inst_funct;
  wire[4:0] Queue_io_deq_bits_inst_rs2;
  wire[4:0] Queue_io_deq_bits_inst_rs1;
  wire Queue_io_deq_bits_inst_xd;
  wire Queue_io_deq_bits_inst_xs1;
  wire Queue_io_deq_bits_inst_xs2;
  wire[4:0] Queue_io_deq_bits_inst_rd;
  wire[6:0] Queue_io_deq_bits_inst_opcode;
  wire[63:0] Queue_io_deq_bits_rs1;
  wire[63:0] Queue_io_deq_bits_rs2;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = cmdReadys_0 <= 1'h1;
  assign cmdReadys_0 = io_out_0_ready & T3;
  assign T3 = 7'hb == Queue_io_deq_bits_inst_opcode;
  assign io_busy = Queue_io_deq_valid;
  assign io_out_0_bits_rs2 = Queue_io_deq_bits_rs2;
  assign io_out_0_bits_rs1 = Queue_io_deq_bits_rs1;
  assign io_out_0_bits_inst_opcode = Queue_io_deq_bits_inst_opcode;
  assign io_out_0_bits_inst_rd = Queue_io_deq_bits_inst_rd;
  assign io_out_0_bits_inst_xs2 = Queue_io_deq_bits_inst_xs2;
  assign io_out_0_bits_inst_xs1 = Queue_io_deq_bits_inst_xs1;
  assign io_out_0_bits_inst_xd = Queue_io_deq_bits_inst_xd;
  assign io_out_0_bits_inst_rs1 = Queue_io_deq_bits_inst_rs1;
  assign io_out_0_bits_inst_rs2 = Queue_io_deq_bits_inst_rs2;
  assign io_out_0_bits_inst_funct = Queue_io_deq_bits_inst_funct;
  assign io_out_0_valid = T4;
  assign T4 = Queue_io_deq_valid & T3;
  assign io_in_ready = Queue_io_enq_ready;
  Queue_10 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_in_valid ),
       .io_enq_bits_inst_funct( io_in_bits_inst_funct ),
       .io_enq_bits_inst_rs2( io_in_bits_inst_rs2 ),
       .io_enq_bits_inst_rs1( io_in_bits_inst_rs1 ),
       .io_enq_bits_inst_xd( io_in_bits_inst_xd ),
       .io_enq_bits_inst_xs1( io_in_bits_inst_xs1 ),
       .io_enq_bits_inst_xs2( io_in_bits_inst_xs2 ),
       .io_enq_bits_inst_rd( io_in_bits_inst_rd ),
       .io_enq_bits_inst_opcode( io_in_bits_inst_opcode ),
       .io_enq_bits_rs1( io_in_bits_rs1 ),
       .io_enq_bits_rs2( io_in_bits_rs2 ),
       .io_deq_ready( cmdReadys_0 ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_inst_funct( Queue_io_deq_bits_inst_funct ),
       .io_deq_bits_inst_rs2( Queue_io_deq_bits_inst_rs2 ),
       .io_deq_bits_inst_rs1( Queue_io_deq_bits_inst_rs1 ),
       .io_deq_bits_inst_xd( Queue_io_deq_bits_inst_xd ),
       .io_deq_bits_inst_xs1( Queue_io_deq_bits_inst_xs1 ),
       .io_deq_bits_inst_xs2( Queue_io_deq_bits_inst_xs2 ),
       .io_deq_bits_inst_rd( Queue_io_deq_bits_inst_rd ),
       .io_deq_bits_inst_opcode( Queue_io_deq_bits_inst_opcode ),
       .io_deq_bits_rs1( Queue_io_deq_bits_rs1 ),
       .io_deq_bits_rs2( Queue_io_deq_bits_rs2 )
       //.io_count(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Custom opcode matched for more than one accelerator");
    $finish;
  end
// synthesis translate_on
`endif
  end
endmodule

// Yangyi: RTL adder
module adder_Accel
(
  clk,
  rst,
  cmd,
  cmd_vld,
  cmd_rdy,
  resp,
  resp_vld,
  resp_rdy,      
);

//  initial begin
//    $display("adder_Accel");
//  end

  // check if can remove the "wire"s
  input              clk;
  input              rst;
  input      [159:0] cmd;
  input              cmd_vld;
  output reg         cmd_rdy;
  output     [73:0]  resp;
  output reg         resp_vld;
  input              resp_rdy;
  
  // Spread The cmd Wires
  wire [6:0]  cmd_inst_funct;  
  wire [4:0]  cmd_inst_rs2;    
  wire [4:0]  cmd_inst_rs1;    
  wire        cmd_inst_xd;     
  wire        cmd_inst_xs1;    
  wire        cmd_inst_xs2;    
  wire [4:0]  cmd_inst_rd;     
  wire [6:0]  cmd_inst_opcode; 
  wire [63:0] cmd_rs1_data;         
  wire [63:0] cmd_rs2_data;         
  
  assign cmd_inst_funct  = cmd[6:0];
  assign cmd_inst_rs2    = cmd[11:7];
  assign cmd_inst_rs1    = cmd[16:12];
  assign cmd_inst_xd     = cmd[17];
  assign cmd_inst_xs1    = cmd[18];
  assign cmd_inst_xs2    = cmd[19];
  assign cmd_inst_rd     = cmd[24:20];
  assign cmd_inst_opcode = cmd[31:25];
  assign cmd_rs1_data    = cmd[95:32];
  assign cmd_rs2_data    = cmd[159:96];
  
  // Generate resp Wires
  wire [63:0] resp_data;
  wire [4:0]  resp_rd;
  wire        SampleAccel_io_mem_req_valid;
  wire        SampleAccel_io_autl_acquire_valid;
  wire        ClientTileLinkIOArbiter_io_in_1_acquire_ready;
  wire        SampleAccel_io_interrupt;
  wire        SampleAccel_io_busy;
  
  assign resp = 
           {
           resp_data, 
           resp_rd, 
           SampleAccel_io_mem_req_valid, 
           SampleAccel_io_autl_acquire_valid, 
           ClientTileLinkIOArbiter_io_in_1_acquire_ready,
           SampleAccel_io_interrupt,
           SampleAccel_io_busy
           };

  // ---Datapath---
  // Add
  parameter data_nbits = 64;
  
  wire [data_nbits-1:0] adder_out;
  
  yh326_Adder#(data_nbits) adder
  (
    .in0 (cmd_rs1_data),
    .in1 (cmd_rs2_data),
    .out (adder_out)
  );
  
  yh326_Reg#(data_nbits) d_reg
  (
    .clk (clk),
    .q   (resp_data),
    .d   (adder_out)
  );
  
  // rd transition
  parameter rd_nbits = 5;
  
  yh326_Reg#(rd_nbits) rd_reg
  (
    .clk (clk),
    .q   (resp_rd),
    .d   (cmd_inst_rd)
  );
  
  // Assign Values To The 5 Unused resp Ports
  assign SampleAccel_io_mem_req_valid = 1'b0;
  assign SampleAccel_io_autl_acquire_valid = 1'b0;
  assign ClientTileLinkIOArbiter_io_in_1_acquire_ready = 1'b0;
  assign SampleAccel_io_interrupt = 1'b0;
  assign SampleAccel_io_busy = 1'b0;

  // ---Control Path---
  // States Definition
  parameter STATE_IDLE = 2'd0;
  parameter STATE_DONE = 2'd1;

  // State Advancement
  reg [1:0]  state_reg;
  reg [1:0]  next_state;

  always @ (posedge clk) begin
    if (rst) begin
      state_reg <= STATE_IDLE;
    end else begin
      state_reg <= next_state;
    end
  end

  // State Advancement Calculations
  wire cmd_go;
  wire resp_go;

  assign cmd_go  = cmd_vld  && cmd_rdy;
  assign resp_go = resp_vld && resp_rdy; 

  always @ (*) begin
    case ( state_reg )
      STATE_IDLE: 
        begin
          if (cmd_go) begin
            next_state = STATE_DONE;
          end else begin
            next_state = state_reg;
          end
        end
      STATE_DONE: 
        begin
          if (resp_go) begin
            next_state = STATE_IDLE;
          end else begin
            next_state = state_reg;
          end
        end
    endcase
  end

  // State Outputs
  always @ (*) begin
    case ( state_reg )
      STATE_IDLE:
        begin
        cmd_rdy  = 1'b1;
        resp_vld = 1'b0;
        end
      STATE_DONE:
        begin
        cmd_rdy  = 1'b0;
        resp_vld = 1'b1;
        end
    endcase
  end
  /*
  task as
  (
    input as_cmd_rdy;
    input as_resp_vld
  );
  begin
    cmd_rdy  = as_cmd_rdy;
    resp_vld = as_resp_vld;
  end
  endtask
  
  always @ (*) begin
    case ( state_reg )
      //              cmd_rdy, resp_vld
      STATE_IDLE:  as(      1,        0);
      STATE_DONE:  as(      0,        1);
    endcase
  end
  */
endmodule

module yh326_Adder
#(
  parameter p_nbits = 1
)(
  in0,
  in1,
  //cin,
  out,
  //cout
);

  input  [p_nbits-1:0] in0;
  input  [p_nbits-1:0] in1;
  //input                cin;
  output [p_nbits-1:0] out;
  //output               cout;

  //assign {cout,out} = in0 + in1 + cin;
  assign out = in0 + in1;

endmodule

module yh326_Reg
#(
  parameter p_nbits = 1
)(
  clk, // Clock input
  q,   // Data output
  d    // Data input
);

  input                    clk;
  output reg [p_nbits-1:0] q;
  input      [p_nbits-1:0] d;

  always @( posedge clk ) begin
    q <= d;
  end

endmodule

//gai: gcd accelerator gererated by vivado HLS

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC
// Version: 2015.3
// Copyright (C) 2015 Xilinx Inc. All rights reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="gcd,hls_ip_2015_3,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xc7z020clg484-2,HLS_INPUT_CLOCK=5.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=3.950000,HLS_SYN_LAT=-1,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=137,HLS_SYN_LUT=430}" *)

module gcd (
        ap_clk,
        ap_rst,
        io_cmd_V,
        io_cmd_V_ap_vld,
        io_cmd_V_ap_ack,
        io_resp_V,
        io_resp_V_ap_vld,
        io_resp_V_ap_ack
);

parameter    ap_const_logic_1 = 1'b1;
parameter    ap_const_logic_0 = 1'b0;
parameter    ap_ST_st1_fsm_0 = 3'b1;
parameter    ap_ST_st2_fsm_1 = 3'b10;
parameter    ap_ST_st3_fsm_2 = 3'b100;
parameter    ap_const_lv32_0 = 32'b00000000000000000000000000000000;
parameter    ap_const_lv1_1 = 1'b1;
parameter    ap_const_lv32_1 = 32'b1;
parameter    ap_const_lv1_0 = 1'b0;
parameter    ap_const_lv32_2 = 32'b10;
parameter    ap_const_lv32_14 = 32'b10100;
parameter    ap_const_lv32_18 = 32'b11000;
parameter    ap_const_lv32_20 = 32'b100000;
parameter    ap_const_lv32_5F = 32'b1011111;
parameter    ap_const_lv32_60 = 32'b1100000;
parameter    ap_const_lv32_9F = 32'b10011111;
parameter    ap_const_lv5_0 = 5'b00000;
parameter    ap_true = 1'b1;

input   ap_clk;
input   ap_rst;
input  [159:0] io_cmd_V;
input   io_cmd_V_ap_vld;
output   io_cmd_V_ap_ack;
output  [73:0] io_resp_V;
output   io_resp_V_ap_vld;
input   io_resp_V_ap_ack;

reg io_cmd_V_ap_ack;
reg io_resp_V_ap_vld;
reg   [4:0] tmp_rd_V_reg_166;
(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm = 3'b1;
reg    ap_sig_cseq_ST_st1_fsm_0;
reg    ap_sig_bdd_24;
wire   [63:0] a_V_2_fu_140_p3;
reg    ap_sig_cseq_ST_st2_fsm_1;
reg    ap_sig_bdd_41;
wire   [0:0] tmp_fu_116_p2;
wire   [63:0] b_V_2_fu_148_p3;
reg   [63:0] tmp_data_V_reg_67;
reg   [63:0] p_1_reg_77;
reg    ap_sig_cseq_ST_st3_fsm_2;
reg    ap_sig_bdd_60;
reg    ap_reg_ioackin_io_resp_V_ap_ack = 1'b0;
reg    ap_sig_ioackin_io_resp_V_ap_ack;
wire   [0:0] tmp_2_fu_122_p2;
wire   [63:0] a_V_1_fu_128_p2;
wire   [63:0] b_V_1_fu_134_p2;
reg   [2:0] ap_NS_fsm;




/// the current state (ap_CS_fsm) of the state machine. ///
always @ (posedge ap_clk) begin : ap_ret_ap_CS_fsm
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_st1_fsm_0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

/// ap_reg_ioackin_io_resp_V_ap_ack assign process. ///
always @ (posedge ap_clk) begin : ap_ret_ap_reg_ioackin_io_resp_V_ap_ack
    if (ap_rst == 1'b1) begin
        ap_reg_ioackin_io_resp_V_ap_ack <= ap_const_logic_0;
    end else begin
        if ((ap_const_logic_1 == ap_sig_cseq_ST_st3_fsm_2)) begin
            if (~(ap_const_logic_0 == ap_sig_ioackin_io_resp_V_ap_ack)) begin
                ap_reg_ioackin_io_resp_V_ap_ack <= ap_const_logic_0;
            end else if ((ap_const_logic_1 == io_resp_V_ap_ack)) begin
                ap_reg_ioackin_io_resp_V_ap_ack <= ap_const_logic_1;
            end
        end
    end
end

/// assign process. ///
always @ (posedge ap_clk) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st2_fsm_1) & (tmp_fu_116_p2 == ap_const_lv1_0))) begin
        p_1_reg_77 <= b_V_2_fu_148_p3;
    end else if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_ap_vld == ap_const_logic_0))) begin
        p_1_reg_77 <= {{io_cmd_V[ap_const_lv32_9F : ap_const_lv32_60]}};
    end
end

/// assign process. ///
always @ (posedge ap_clk) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st2_fsm_1) & (tmp_fu_116_p2 == ap_const_lv1_0))) begin
        tmp_data_V_reg_67 <= a_V_2_fu_140_p3;
    end else if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_ap_vld == ap_const_logic_0))) begin
        tmp_data_V_reg_67 <= {{io_cmd_V[ap_const_lv32_5F : ap_const_lv32_20]}};
    end
end

/// assign process. ///
always @ (posedge ap_clk) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_ap_vld == ap_const_logic_0))) begin
        tmp_rd_V_reg_166 <= {{io_cmd_V[ap_const_lv32_18 : ap_const_lv32_14]}};
    end
end

/// ap_sig_cseq_ST_st1_fsm_0 assign process. ///
always @ (ap_sig_bdd_24) begin
    if (ap_sig_bdd_24) begin
        ap_sig_cseq_ST_st1_fsm_0 = ap_const_logic_1;
    end else begin
        ap_sig_cseq_ST_st1_fsm_0 = ap_const_logic_0;
    end
end

/// ap_sig_cseq_ST_st2_fsm_1 assign process. ///
always @ (ap_sig_bdd_41) begin
    if (ap_sig_bdd_41) begin
        ap_sig_cseq_ST_st2_fsm_1 = ap_const_logic_1;
    end else begin
        ap_sig_cseq_ST_st2_fsm_1 = ap_const_logic_0;
    end
end

/// ap_sig_cseq_ST_st3_fsm_2 assign process. ///
always @ (ap_sig_bdd_60) begin
    if (ap_sig_bdd_60) begin
        ap_sig_cseq_ST_st3_fsm_2 = ap_const_logic_1;
    end else begin
        ap_sig_cseq_ST_st3_fsm_2 = ap_const_logic_0;
    end
end

/// ap_sig_ioackin_io_resp_V_ap_ack assign process. ///
always @ (io_resp_V_ap_ack or ap_reg_ioackin_io_resp_V_ap_ack) begin
    if ((ap_const_logic_0 == ap_reg_ioackin_io_resp_V_ap_ack)) begin
        ap_sig_ioackin_io_resp_V_ap_ack = io_resp_V_ap_ack;
    end else begin
        ap_sig_ioackin_io_resp_V_ap_ack = ap_const_logic_1;
    end
end

/// io_cmd_V_ap_ack assign process. ///
always @ (io_cmd_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_ap_vld == ap_const_logic_0))) begin
        io_cmd_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_ap_ack = ap_const_logic_0;
    end
end

/// io_resp_V_ap_vld assign process. ///
always @ (ap_sig_cseq_ST_st3_fsm_2 or ap_reg_ioackin_io_resp_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st3_fsm_2) & (ap_const_logic_0 == ap_reg_ioackin_io_resp_V_ap_ack))) begin
        io_resp_V_ap_vld = ap_const_logic_1;
    end else begin
        io_resp_V_ap_vld = ap_const_logic_0;
    end
end
/// the next state (ap_NS_fsm) of the state machine. ///
always @ (io_cmd_V_ap_vld or ap_CS_fsm or tmp_fu_116_p2 or ap_sig_ioackin_io_resp_V_ap_ack) begin
    case (ap_CS_fsm)
        ap_ST_st1_fsm_0 : 
        begin
            if (~(io_cmd_V_ap_vld == ap_const_logic_0)) begin
                ap_NS_fsm = ap_ST_st2_fsm_1;
            end else begin
                ap_NS_fsm = ap_ST_st1_fsm_0;
            end
        end
        ap_ST_st2_fsm_1 : 
        begin
            if ((tmp_fu_116_p2 == ap_const_lv1_0)) begin
                ap_NS_fsm = ap_ST_st2_fsm_1;
            end else begin
                ap_NS_fsm = ap_ST_st3_fsm_2;
            end
        end
        ap_ST_st3_fsm_2 : 
        begin
            if (~(ap_const_logic_0 == ap_sig_ioackin_io_resp_V_ap_ack)) begin
                ap_NS_fsm = ap_ST_st1_fsm_0;
            end else begin
                ap_NS_fsm = ap_ST_st3_fsm_2;
            end
        end
        default : 
        begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign a_V_1_fu_128_p2 = (tmp_data_V_reg_67 - p_1_reg_77);
assign a_V_2_fu_140_p3 = ((tmp_2_fu_122_p2[0:0] === 1'b1) ? a_V_1_fu_128_p2 : tmp_data_V_reg_67);

/// ap_sig_bdd_24 assign process. ///
always @ (ap_CS_fsm) begin
    ap_sig_bdd_24 = (ap_CS_fsm[ap_const_lv32_0] == ap_const_lv1_1);
end

/// ap_sig_bdd_41 assign process. ///
always @ (ap_CS_fsm) begin
    ap_sig_bdd_41 = (ap_const_lv1_1 == ap_CS_fsm[ap_const_lv32_1]);
end

/// ap_sig_bdd_60 assign process. ///
always @ (ap_CS_fsm) begin
    ap_sig_bdd_60 = (ap_const_lv1_1 == ap_CS_fsm[ap_const_lv32_2]);
end
assign b_V_1_fu_134_p2 = (p_1_reg_77 - tmp_data_V_reg_67);
assign b_V_2_fu_148_p3 = ((tmp_2_fu_122_p2[0:0] === 1'b1) ? p_1_reg_77 : b_V_1_fu_134_p2);
assign io_resp_V = {{{tmp_data_V_reg_67}, {tmp_rd_V_reg_166}}, {ap_const_lv5_0}};
assign tmp_2_fu_122_p2 = (tmp_data_V_reg_67 > p_1_reg_77? 1'b1: 1'b0);
assign tmp_fu_116_p2 = (tmp_data_V_reg_67 == p_1_reg_77? 1'b1: 1'b0);


endmodule //gcd

// ==============================================================
// RTL generated by Vivado(TM) HLS - High-Level Synthesis from C, C++ and SystemC
// Version: 2015.3
// Copyright (C) 2015 Xilinx Inc. All rights reserved.
// 
// ===========================================================

module add (
        ap_clk,
        ap_rst,
        io_cmd_V_inst_funct_V,
        io_cmd_V_inst_funct_V_ap_vld,
        io_cmd_V_inst_funct_V_ap_ack,
        io_cmd_V_inst_rs2_V,
        io_cmd_V_inst_rs2_V_ap_vld,
        io_cmd_V_inst_rs2_V_ap_ack,
        io_cmd_V_inst_rs1_V,
        io_cmd_V_inst_rs1_V_ap_vld,
        io_cmd_V_inst_rs1_V_ap_ack,
        io_cmd_V_inst_xd_V,
        io_cmd_V_inst_xd_V_ap_vld,
        io_cmd_V_inst_xd_V_ap_ack,
        io_cmd_V_inst_xs1_V,
        io_cmd_V_inst_xs1_V_ap_vld,
        io_cmd_V_inst_xs1_V_ap_ack,
        io_cmd_V_inst_xs2_V,
        io_cmd_V_inst_xs2_V_ap_vld,
        io_cmd_V_inst_xs2_V_ap_ack,
        io_cmd_V_inst_rd_V,
        io_cmd_V_inst_rd_V_ap_vld,
        io_cmd_V_inst_rd_V_ap_ack,
        io_cmd_V_inst_opcode_V,
        io_cmd_V_inst_opcode_V_ap_vld,
        io_cmd_V_inst_opcode_V_ap_ack,
        io_cmd_V_rs1_V,
        io_cmd_V_rs1_V_ap_vld,
        io_cmd_V_rs1_V_ap_ack,
        io_cmd_V_rs2_V,
        io_cmd_V_rs2_V_ap_vld,
        io_cmd_V_rs2_V_ap_ack,
        io_resp_V_rd_V,
        io_resp_V_rd_V_ap_vld,
        io_resp_V_rd_V_ap_ack,
        io_resp_V_data_V,
        io_resp_V_data_V_ap_vld,
        io_resp_V_data_V_ap_ack,
        io_mem_req_ready,
        io_mem_req_valid,
        io_busy,
        io_interrupt,
        io_autl_acquire_ready,
        io_autl_acquire_valid
);

parameter    ap_const_logic_1 = 1'b1;
parameter    ap_const_logic_0 = 1'b0;
parameter    ap_ST_st1_fsm_0 = 1'b1;
parameter    ap_const_lv32_0 = 32'b00000000000000000000000000000000;
parameter    ap_const_lv1_1 = 1'b1;
parameter    ap_true = 1'b1;

input   ap_clk;
input   ap_rst;
input  [6:0] io_cmd_V_inst_funct_V;
input   io_cmd_V_inst_funct_V_ap_vld;
output   io_cmd_V_inst_funct_V_ap_ack;
input  [4:0] io_cmd_V_inst_rs2_V;
input   io_cmd_V_inst_rs2_V_ap_vld;
output   io_cmd_V_inst_rs2_V_ap_ack;
input  [4:0] io_cmd_V_inst_rs1_V;
input   io_cmd_V_inst_rs1_V_ap_vld;
output   io_cmd_V_inst_rs1_V_ap_ack;
input  [0:0] io_cmd_V_inst_xd_V;
input   io_cmd_V_inst_xd_V_ap_vld;
output   io_cmd_V_inst_xd_V_ap_ack;
input  [0:0] io_cmd_V_inst_xs1_V;
input   io_cmd_V_inst_xs1_V_ap_vld;
output   io_cmd_V_inst_xs1_V_ap_ack;
input  [0:0] io_cmd_V_inst_xs2_V;
input   io_cmd_V_inst_xs2_V_ap_vld;
output   io_cmd_V_inst_xs2_V_ap_ack;
input  [4:0] io_cmd_V_inst_rd_V;
input   io_cmd_V_inst_rd_V_ap_vld;
output   io_cmd_V_inst_rd_V_ap_ack;
input  [6:0] io_cmd_V_inst_opcode_V;
input   io_cmd_V_inst_opcode_V_ap_vld;
output   io_cmd_V_inst_opcode_V_ap_ack;
input  [63:0] io_cmd_V_rs1_V;
input   io_cmd_V_rs1_V_ap_vld;
output   io_cmd_V_rs1_V_ap_ack;
input  [63:0] io_cmd_V_rs2_V;
input   io_cmd_V_rs2_V_ap_vld;
output   io_cmd_V_rs2_V_ap_ack;
output  [4:0] io_resp_V_rd_V;
output   io_resp_V_rd_V_ap_vld;
input   io_resp_V_rd_V_ap_ack;
output  [63:0] io_resp_V_data_V;
output   io_resp_V_data_V_ap_vld;
input   io_resp_V_data_V_ap_ack;

output io_busy;
output io_interrupt;
output io_autl_acquire_ready;
output io_autl_acquire_valid;
output io_mem_req_valid;
input io_mem_req_ready;

assign io_autl_grant_ready = 1'h0;
assign io_autl_acquire_valid = 1'h0;
assign io_interrupt = 1'h0;
assign io_busy = 1'h0;
assign io_mem_req_valid = 1'h0; 

reg io_cmd_V_inst_funct_V_ap_ack;
reg io_cmd_V_inst_rs2_V_ap_ack;
reg io_cmd_V_inst_rs1_V_ap_ack;
reg io_cmd_V_inst_xd_V_ap_ack;
reg io_cmd_V_inst_xs1_V_ap_ack;
reg io_cmd_V_inst_xs2_V_ap_ack;
reg io_cmd_V_inst_rd_V_ap_ack;
reg io_cmd_V_inst_opcode_V_ap_ack;
reg io_cmd_V_rs1_V_ap_ack;
reg io_cmd_V_rs2_V_ap_ack;
reg io_resp_V_rd_V_ap_vld;
reg io_resp_V_data_V_ap_vld;
(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm = 1'b1;
reg    ap_sig_cseq_ST_st1_fsm_0;
reg    ap_sig_bdd_61;
reg    ap_sig_ioackin_io_resp_V_rd_V_ap_ack;
reg    ap_reg_ioackin_io_resp_V_rd_V_ap_ack = 1'b0;
reg    ap_reg_ioackin_io_resp_V_data_V_ap_ack = 1'b0;
reg   [0:0] ap_NS_fsm;
reg    ap_sig_bdd_133;
reg    ap_sig_bdd_135;

/// the current state (ap_CS_fsm) of the state machine. ///
always @ (posedge ap_clk) begin : ap_ret_ap_CS_fsm
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_st1_fsm_0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

/// ap_reg_ioackin_io_resp_V_data_V_ap_ack assign process. ///
always @ (posedge ap_clk) begin : ap_ret_ap_reg_ioackin_io_resp_V_data_V_ap_ack
    if (ap_rst == 1'b1) begin
        ap_reg_ioackin_io_resp_V_data_V_ap_ack <= ap_const_logic_0;
    end else begin
        if ((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0)) begin
            if (~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack))) begin
                ap_reg_ioackin_io_resp_V_data_V_ap_ack <= ap_const_logic_0;
            end else if (ap_sig_bdd_133) begin
                ap_reg_ioackin_io_resp_V_data_V_ap_ack <= ap_const_logic_1;
            end
        end
    end
end

/// ap_reg_ioackin_io_resp_V_rd_V_ap_ack assign process. ///
always @ (posedge ap_clk) begin : ap_ret_ap_reg_ioackin_io_resp_V_rd_V_ap_ack
    if (ap_rst == 1'b1) begin
        ap_reg_ioackin_io_resp_V_rd_V_ap_ack <= ap_const_logic_0;
    end else begin
        if ((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0)) begin
            if (~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack))) begin
                ap_reg_ioackin_io_resp_V_rd_V_ap_ack <= ap_const_logic_0;
            end else if (ap_sig_bdd_135) begin
                ap_reg_ioackin_io_resp_V_rd_V_ap_ack <= ap_const_logic_1;
            end
        end
    end
end

/// ap_sig_cseq_ST_st1_fsm_0 assign process. ///
always @ (ap_sig_bdd_61) begin
    if (ap_sig_bdd_61) begin
        ap_sig_cseq_ST_st1_fsm_0 = ap_const_logic_1;
    end else begin
        ap_sig_cseq_ST_st1_fsm_0 = ap_const_logic_0;
    end
end

/// ap_sig_ioackin_io_resp_V_rd_V_ap_ack assign process. ///
always @ (io_resp_V_rd_V_ap_ack or ap_reg_ioackin_io_resp_V_rd_V_ap_ack) begin
    if ((ap_const_logic_0 == ap_reg_ioackin_io_resp_V_rd_V_ap_ack)) begin
        ap_sig_ioackin_io_resp_V_rd_V_ap_ack = io_resp_V_rd_V_ap_ack;
    end else begin
        ap_sig_ioackin_io_resp_V_rd_V_ap_ack = ap_const_logic_1;
    end
end

/// io_cmd_V_inst_funct_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_funct_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_funct_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_opcode_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_opcode_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_opcode_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_rd_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_rd_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_rd_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_rs1_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_rs1_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_rs1_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_rs2_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_rs2_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_rs2_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_xd_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_xd_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_xd_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_xs1_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_xs1_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_xs1_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_inst_xs2_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_inst_xs2_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_inst_xs2_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_rs1_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_rs1_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_rs1_V_ap_ack = ap_const_logic_0;
    end
end

/// io_cmd_V_rs2_V_ap_ack assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~((io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) | (ap_const_logic_0 == ap_sig_ioackin_io_resp_V_rd_V_ap_ack)))) begin
        io_cmd_V_rs2_V_ap_ack = ap_const_logic_1;
    end else begin
        io_cmd_V_rs2_V_ap_ack = ap_const_logic_0;
    end
end

/// io_resp_V_data_V_ap_vld assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_reg_ioackin_io_resp_V_data_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) & (ap_const_logic_0 == ap_reg_ioackin_io_resp_V_data_V_ap_ack))) begin
        io_resp_V_data_V_ap_vld = ap_const_logic_1;
    end else begin
        io_resp_V_data_V_ap_vld = ap_const_logic_0;
    end
end

/// io_resp_V_rd_V_ap_vld assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_sig_cseq_ST_st1_fsm_0 or ap_reg_ioackin_io_resp_V_rd_V_ap_ack) begin
    if (((ap_const_logic_1 == ap_sig_cseq_ST_st1_fsm_0) & ~(io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) & (ap_const_logic_0 == ap_reg_ioackin_io_resp_V_rd_V_ap_ack))) begin
        io_resp_V_rd_V_ap_vld = ap_const_logic_1;
    end else begin
        io_resp_V_rd_V_ap_vld = ap_const_logic_0;
    end
end
/// the next state (ap_NS_fsm) of the state machine. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or ap_CS_fsm or ap_sig_ioackin_io_resp_V_rd_V_ap_ack) begin
    case (ap_CS_fsm)
        ap_ST_st1_fsm_0 : 
        begin
            ap_NS_fsm = ap_ST_st1_fsm_0;
        end
        default : 
        begin
            ap_NS_fsm = 'bx;
        end
    endcase
end


/// ap_sig_bdd_133 assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or io_resp_V_data_V_ap_ack) begin
    ap_sig_bdd_133 = (~(io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) & (ap_const_logic_1 == io_resp_V_data_V_ap_ack));
end

/// ap_sig_bdd_135 assign process. ///
always @ (io_cmd_V_inst_funct_V_ap_vld or io_resp_V_rd_V_ap_ack) begin
    ap_sig_bdd_135 = (~(io_cmd_V_inst_funct_V_ap_vld == ap_const_logic_0) & (ap_const_logic_1 == io_resp_V_rd_V_ap_ack));
end

/// ap_sig_bdd_61 assign process. ///
always @ (ap_CS_fsm) begin
    ap_sig_bdd_61 = (ap_CS_fsm[ap_const_lv32_0] == ap_const_lv1_1);
end
assign io_resp_V_data_V = (io_cmd_V_rs2_V + io_cmd_V_rs1_V);
assign io_resp_V_rd_V = io_cmd_V_inst_rd_V;


endmodule //add


/*
module SampleAccel(input clk, input reset,
    output io_cmd_ready,
    input  io_cmd_valid,
    input [6:0] io_cmd_bits_inst_funct,
    input [4:0] io_cmd_bits_inst_rs2,
    input [4:0] io_cmd_bits_inst_rs1,
    input  io_cmd_bits_inst_xd,
    input  io_cmd_bits_inst_xs1,
    input  io_cmd_bits_inst_xs2,
    input [4:0] io_cmd_bits_inst_rd,
    input [6:0] io_cmd_bits_inst_opcode,
    input [63:0] io_cmd_bits_rs1,
    input [63:0] io_cmd_bits_rs2,
    input  io_resp_ready,
    output io_resp_valid,
    output[4:0] io_resp_bits_rd,
    output[63:0] io_resp_bits_data,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    //output[39:0] io_mem_req_bits_addr
    //output[9:0] io_mem_req_bits_tag
    //output[4:0] io_mem_req_bits_cmd
    //output[2:0] io_mem_req_bits_typ
    //output io_mem_req_bits_kill
    output io_mem_req_bits_phys,
    //output[63:0] io_mem_req_bits_data
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [9:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    //input  io_mem_replay_next_valid
    //input [9:0] io_mem_replay_next_bits
    //input  io_mem_xcpt_ma_ld
    //input  io_mem_xcpt_ma_st
    //input  io_mem_xcpt_pf_ld
    //input  io_mem_xcpt_pf_st
    //output io_mem_invalidate_lr
    //input  io_mem_ordered
    output io_busy,
    input  io_s,
    output io_interrupt,
    input  io_autl_acquire_ready,
    output io_autl_acquire_valid,
    //output[25:0] io_autl_acquire_bits_addr_block
    //output[5:0] io_autl_acquire_bits_client_xact_id
    //output[1:0] io_autl_acquire_bits_addr_beat
    //output io_autl_acquire_bits_is_builtin_type
    //output[2:0] io_autl_acquire_bits_a_type
    //output[16:0] io_autl_acquire_bits_union
    //output[127:0] io_autl_acquire_bits_data
    output io_autl_grant_ready,
    input  io_autl_grant_valid,
    input [1:0] io_autl_grant_bits_addr_beat,
    input [5:0] io_autl_grant_bits_client_xact_id,
    input [3:0] io_autl_grant_bits_manager_xact_id,
    input  io_autl_grant_bits_is_builtin_type,
    input [3:0] io_autl_grant_bits_g_type,
    input [127:0] io_autl_grant_bits_data,
    //input  io_fpu_req_ready
    //output io_fpu_req_valid
    //output[4:0] io_fpu_req_bits_cmd
    //output io_fpu_req_bits_ldst
    //output io_fpu_req_bits_wen
    //output io_fpu_req_bits_ren1
    //output io_fpu_req_bits_ren2
    //output io_fpu_req_bits_ren3
    //output io_fpu_req_bits_swap12
    //output io_fpu_req_bits_swap23
    //output io_fpu_req_bits_single
    //output io_fpu_req_bits_fromint
    //output io_fpu_req_bits_toint
    //output io_fpu_req_bits_fastpipe
    //output io_fpu_req_bits_fma
    //output io_fpu_req_bits_div
    //output io_fpu_req_bits_sqrt
    //output io_fpu_req_bits_round
    //output io_fpu_req_bits_wflags
    //output[2:0] io_fpu_req_bits_rm
    //output[1:0] io_fpu_req_bits_typ
    //output[64:0] io_fpu_req_bits_in1
    //output[64:0] io_fpu_req_bits_in2
    //output[64:0] io_fpu_req_bits_in3
    //output io_fpu_resp_ready
    //input  io_fpu_resp_valid
    //input [64:0] io_fpu_resp_bits_data
    //input [4:0] io_fpu_resp_bits_exc
    input  io_exception,
    //input [11:0] io_csr_waddr
    //input [63:0] io_csr_wdata
    //input  io_csr_wen
    input  io_host_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg  state;
  wire T62;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] T33;
  reg [63:0] rs2_reg;
  wire[63:0] T63;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  reg [63:0] rs1_reg;
  wire[63:0] T64;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[4:0] T45;
  wire[4:0] T46;
  wire[4:0] T47;
  wire[4:0] T48;
  reg [4:0] rd_reg;
  wire[4:0] T65;
  wire[4:0] T49;
  wire[4:0] T50;
  wire[4:0] T51;
  wire[4:0] T52;
  wire[4:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    rs2_reg = {2{$random}};
    rs1_reg = {2{$random}};
    rd_reg = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_fpu_resp_ready = {1{$random}};
//  assign io_fpu_req_bits_in3 = {3{$random}};
//  assign io_fpu_req_bits_in2 = {3{$random}};
//  assign io_fpu_req_bits_in1 = {3{$random}};
//  assign io_fpu_req_bits_typ = {1{$random}};
//  assign io_fpu_req_bits_rm = {1{$random}};
//  assign io_fpu_req_bits_wflags = {1{$random}};
//  assign io_fpu_req_bits_round = {1{$random}};
//  assign io_fpu_req_bits_sqrt = {1{$random}};
//  assign io_fpu_req_bits_div = {1{$random}};
//  assign io_fpu_req_bits_fma = {1{$random}};
//  assign io_fpu_req_bits_fastpipe = {1{$random}};
//  assign io_fpu_req_bits_toint = {1{$random}};
//  assign io_fpu_req_bits_fromint = {1{$random}};
//  assign io_fpu_req_bits_single = {1{$random}};
//  assign io_fpu_req_bits_swap23 = {1{$random}};
//  assign io_fpu_req_bits_swap12 = {1{$random}};
//  assign io_fpu_req_bits_ren3 = {1{$random}};
//  assign io_fpu_req_bits_ren2 = {1{$random}};
//  assign io_fpu_req_bits_ren1 = {1{$random}};
//  assign io_fpu_req_bits_wen = {1{$random}};
//  assign io_fpu_req_bits_ldst = {1{$random}};
//  assign io_fpu_req_bits_cmd = {1{$random}};
//  assign io_fpu_req_valid = {1{$random}};
//  assign io_autl_acquire_bits_data = {4{$random}};
//  assign io_autl_acquire_bits_union = {1{$random}};
//  assign io_autl_acquire_bits_a_type = {1{$random}};
//  assign io_autl_acquire_bits_is_builtin_type = {1{$random}};
//  assign io_autl_acquire_bits_addr_beat = {1{$random}};
//  assign io_autl_acquire_bits_client_xact_id = {1{$random}};
//  assign io_autl_acquire_bits_addr_block = {1{$random}};
//  assign io_mem_invalidate_lr = {1{$random}};
//  assign io_mem_req_bits_data = {2{$random}};
//  assign io_mem_req_bits_kill = {1{$random}};
//  assign io_mem_req_bits_typ = {1{$random}};
//  assign io_mem_req_bits_cmd = {1{$random}};
//  assign io_mem_req_bits_tag = {1{$random}};
//  assign io_mem_req_bits_addr = {2{$random}};
// synthesis translate_on
`endif
  assign io_autl_grant_ready = 1'h0;
  assign io_autl_acquire_valid = 1'h0;
  assign io_interrupt = 1'h0;
  assign io_busy = T0;
  assign T0 = T27 ? 1'h1 : T1;
  assign T1 = T25 ? 1'h1 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h0 : 1'h0;
  assign T4 = T5 & io_cmd_valid;
  assign T5 = state == 1'h0;
  assign T62 = reset ? 1'h0 : T6;
  assign T6 = T11 ? 1'h0 : T7;
  assign T7 = T27 ? 1'h1 : T8;
  assign T8 = T25 ? 1'h0 : T9;
  assign T9 = T23 ? 1'h0 : T10;
  assign T10 = T4 ? 1'h1 : state;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T16 | T13;
  assign T13 = T15 & T14;
  assign T14 = io_resp_ready ^ 1'h1;
  assign T15 = state == 1'h1;
  assign T16 = T19 | T17;
  assign T17 = T18 & io_resp_ready;
  assign T18 = state == 1'h1;
  assign T19 = T4 | T20;
  assign T20 = T22 & T21;
  assign T21 = io_cmd_valid ^ 1'h1;
  assign T22 = state == 1'h0;
  assign T23 = T24 & T20;
  assign T24 = T4 ^ 1'h1;
  assign T25 = T26 & T17;
  assign T26 = T19 ^ 1'h1;
  assign T27 = T28 & T13;
  assign T28 = T16 ^ 1'h1;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_valid = 1'h0;
  assign io_resp_bits_data = T29;
  assign T29 = T27 ? T44 : T30;
  assign T30 = T25 ? T33 : T31;
  assign T31 = T23 ? 64'hf : T32;
  assign T32 = T4 ? 64'hf : 64'hf;
  assign T33 = rs1_reg + rs2_reg;
  assign T63 = reset ? 64'h0 : T34;
  assign T34 = T11 ? rs2_reg : T35;
  assign T35 = T27 ? rs2_reg : T36;
  assign T36 = T25 ? rs2_reg : T37;
  assign T37 = T23 ? io_cmd_bits_rs2 : T38;
  assign T38 = T4 ? io_cmd_bits_rs2 : rs2_reg;
  assign T64 = reset ? 64'h0 : T39;
  assign T39 = T11 ? rs1_reg : T40;
  assign T40 = T27 ? rs1_reg : T41;
  assign T41 = T25 ? rs1_reg : T42;
  assign T42 = T23 ? io_cmd_bits_rs1 : T43;
  assign T43 = T4 ? io_cmd_bits_rs1 : rs1_reg;
  assign T44 = rs1_reg + rs2_reg;
  assign io_resp_bits_rd = T45;
  assign T45 = T27 ? rd_reg : T46;
  assign T46 = T25 ? rd_reg : T47;
  assign T47 = T23 ? 5'h0 : T48;
  assign T48 = T4 ? 5'h0 : 5'h0;
  assign T65 = reset ? 5'h0 : T49;
  assign T49 = T11 ? rd_reg : T50;
  assign T50 = T27 ? rd_reg : T51;
  assign T51 = T25 ? rd_reg : T52;
  assign T52 = T23 ? io_cmd_bits_inst_rd : T53;
  assign T53 = T4 ? io_cmd_bits_inst_rd : rd_reg;
  assign io_resp_valid = T54;
  assign T54 = T27 ? 1'h0 : T55;
  assign T55 = T25 ? 1'h1 : T56;
  assign T56 = T23 ? 1'h0 : T57;
  assign T57 = T4 ? 1'h0 : 1'h0;
  assign io_cmd_ready = T58;
  assign T58 = T27 ? 1'h0 : T59;
  assign T59 = T25 ? 1'h0 : T60;
  assign T60 = T23 ? 1'h1 : T61;
  assign T61 = T4 ? 1'h1 : 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 1'h0;
    end else if(T11) begin
      state <= 1'h0;
    end else if(T27) begin
      state <= 1'h1;
    end else if(T25) begin
      state <= 1'h0;
    end else if(T23) begin
      state <= 1'h0;
    end else if(T4) begin
      state <= 1'h1;
    end
    if(reset) begin
      rs2_reg <= 64'h0;
    end else if(T11) begin
      rs2_reg <= rs2_reg;
    end else if(T27) begin
      rs2_reg <= rs2_reg;
    end else if(T25) begin
      rs2_reg <= rs2_reg;
    end else if(T23) begin
      rs2_reg <= io_cmd_bits_rs2;
    end else if(T4) begin
      rs2_reg <= io_cmd_bits_rs2;
    end
    if(reset) begin
      rs1_reg <= 64'h0;
    end else if(T11) begin
      rs1_reg <= rs1_reg;
    end else if(T27) begin
      rs1_reg <= rs1_reg;
    end else if(T25) begin
      rs1_reg <= rs1_reg;
    end else if(T23) begin
      rs1_reg <= io_cmd_bits_rs1;
    end else if(T4) begin
      rs1_reg <= io_cmd_bits_rs1;
    end
    if(reset) begin
      rd_reg <= 5'h0;
    end else if(T11) begin
      rd_reg <= rd_reg;
    end else if(T27) begin
      rd_reg <= rd_reg;
    end else if(T25) begin
      rd_reg <= rd_reg;
    end else if(T23) begin
      rd_reg <= io_cmd_bits_inst_rd;
    end else if(T4) begin
      rd_reg <= io_cmd_bits_inst_rd;
    end
  end
endmodule
*/


module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [9:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[9:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[63:0] io_deq_bits_data,
    output io_count
);

  wire T33;
  wire[1:0] T0;
  reg  full;
  wire T34;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_flow;
  wire empty;
  wire T3;
  wire T4;
  wire do_deq;
  wire T5;
  wire T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[123:0] T9;
  reg [123:0] ram [0:0];
  wire[123:0] T10;
  wire[123:0] T11;
  wire[123:0] T12;
  wire[68:0] T13;
  wire[64:0] T14;
  wire[3:0] T15;
  wire[54:0] T16;
  wire[14:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[4:0] T24;
  wire[4:0] T25;
  wire[9:0] T26;
  wire[9:0] T27;
  wire[39:0] T28;
  wire[39:0] T29;
  wire T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T33;
  assign T33 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T34 = reset ? 1'h0 : T1;
  assign T1 = T4 ? do_enq : full;
  assign do_enq = T3 & T2;
  assign T2 = do_flow ^ 1'h1;
  assign do_flow = empty & io_deq_ready;
  assign empty = full ^ 1'h1;
  assign T3 = io_enq_ready & io_enq_valid;
  assign T4 = do_enq != do_deq;
  assign do_deq = T6 & T5;
  assign T5 = do_flow ^ 1'h1;
  assign T6 = io_deq_ready & io_deq_valid;
  assign io_deq_bits_data = T7;
  assign T7 = empty ? io_enq_bits_data : T8;
  assign T8 = T9[6'h3f:1'h0];
  assign T9 = ram[1'h0];
  assign T11 = T12;
  assign T12 = {T16, T13};
  assign T13 = {T15, T14};
  assign T14 = {io_enq_bits_phys, io_enq_bits_data};
  assign T15 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T16 = {io_enq_bits_addr, T17};
  assign T17 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T18;
  assign T18 = empty ? io_enq_bits_phys : T19;
  assign T19 = T9[7'h40];
  assign io_deq_bits_kill = T20;
  assign T20 = empty ? io_enq_bits_kill : T21;
  assign T21 = T9[7'h41];
  assign io_deq_bits_typ = T22;
  assign T22 = empty ? io_enq_bits_typ : T23;
  assign T23 = T9[7'h44:7'h42];
  assign io_deq_bits_cmd = T24;
  assign T24 = empty ? io_enq_bits_cmd : T25;
  assign T25 = T9[7'h49:7'h45];
  assign io_deq_bits_tag = T26;
  assign T26 = empty ? io_enq_bits_tag : T27;
  assign T27 = T9[7'h53:7'h4a];
  assign io_deq_bits_addr = T28;
  assign T28 = empty ? io_enq_bits_addr : T29;
  assign T29 = T9[7'h7b:7'h54];
  assign io_deq_valid = T30;
  assign T30 = T31 | io_enq_valid;
  assign T31 = empty ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T4) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T11;
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [9:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[9:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[63:0] io_deq_bits_data,
    output io_count
);

  wire T21;
  wire[1:0] T0;
  reg  full;
  wire T22;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[63:0] T3;
  wire[123:0] T4;
  reg [123:0] ram [0:0];
  wire[123:0] T5;
  wire[123:0] T6;
  wire[123:0] T7;
  wire[68:0] T8;
  wire[64:0] T9;
  wire[3:0] T10;
  wire[54:0] T11;
  wire[14:0] T12;
  wire T13;
  wire T14;
  wire[2:0] T15;
  wire[4:0] T16;
  wire[9:0] T17;
  wire[39:0] T18;
  wire T19;
  wire empty;
  wire T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T21;
  assign T21 = T0[1'h0];
  assign T0 = {full, 1'h0};
  assign T22 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_data = T3;
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_phys, io_enq_bits_data};
  assign T10 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T11 = {io_enq_bits_addr, T12};
  assign T12 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T13;
  assign T13 = T4[7'h40];
  assign io_deq_bits_kill = T14;
  assign T14 = T4[7'h41];
  assign io_deq_bits_typ = T15;
  assign T15 = T4[7'h44:7'h42];
  assign io_deq_bits_cmd = T16;
  assign T16 = T4[7'h49:7'h45];
  assign io_deq_bits_tag = T17;
  assign T17 = T4[7'h53:7'h4a];
  assign io_deq_bits_addr = T18;
  assign T18 = T4[7'h7b:7'h54];
  assign io_deq_valid = T19;
  assign T19 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [39:0] io_in_1_bits_addr,
    input [9:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_kill,
    input  io_in_1_bits_phys,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [9:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_kill,
    input  io_in_0_bits_phys,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[9:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output io_out_bits_kill,
    output io_out_bits_phys,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[63:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire[4:0] T5;
  wire[9:0] T6;
  wire[39:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_phys = T2;
  assign T2 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_kill = T3;
  assign T3 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_bits_typ = T4;
  assign T4 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_cmd = T5;
  assign T5 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T6;
  assign T6 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T7;
  assign T7 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module SimpleHellaCacheIF(input clk, input reset,
    output io_requestor_req_ready,
    input  io_requestor_req_valid,
    input [39:0] io_requestor_req_bits_addr,
    input [9:0] io_requestor_req_bits_tag,
    input [4:0] io_requestor_req_bits_cmd,
    input [2:0] io_requestor_req_bits_typ,
    input  io_requestor_req_bits_kill,
    input  io_requestor_req_bits_phys,
    input [63:0] io_requestor_req_bits_data,
    output io_requestor_resp_valid,
    output[39:0] io_requestor_resp_bits_addr,
    output[9:0] io_requestor_resp_bits_tag,
    output[4:0] io_requestor_resp_bits_cmd,
    output[2:0] io_requestor_resp_bits_typ,
    output[63:0] io_requestor_resp_bits_data,
    output io_requestor_resp_bits_nack,
    output io_requestor_resp_bits_replay,
    output io_requestor_resp_bits_has_data,
    output[63:0] io_requestor_resp_bits_data_word_bypass,
    output[63:0] io_requestor_resp_bits_store_data,
    //output io_requestor_replay_next_valid
    //output[9:0] io_requestor_replay_next_bits
    //output io_requestor_xcpt_ma_ld
    //output io_requestor_xcpt_ma_st
    //output io_requestor_xcpt_pf_ld
    //output io_requestor_xcpt_pf_st
    //input  io_requestor_invalidate_lr
    //output io_requestor_ordered
    input  io_cache_req_ready,
    output io_cache_req_valid,
    output[39:0] io_cache_req_bits_addr,
    output[9:0] io_cache_req_bits_tag,
    output[4:0] io_cache_req_bits_cmd,
    output[2:0] io_cache_req_bits_typ,
    output io_cache_req_bits_kill,
    output io_cache_req_bits_phys,
    output[63:0] io_cache_req_bits_data,
    input  io_cache_resp_valid,
    input [39:0] io_cache_resp_bits_addr,
    input [9:0] io_cache_resp_bits_tag,
    input [4:0] io_cache_resp_bits_cmd,
    input [2:0] io_cache_resp_bits_typ,
    input [63:0] io_cache_resp_bits_data,
    input  io_cache_resp_bits_nack,
    input  io_cache_resp_bits_replay,
    input  io_cache_resp_bits_has_data,
    input [63:0] io_cache_resp_bits_data_word_bypass,
    input [63:0] io_cache_resp_bits_store_data,
    input  io_cache_replay_next_valid,
    input [9:0] io_cache_replay_next_bits,
    input  io_cache_xcpt_ma_ld,
    input  io_cache_xcpt_ma_st,
    input  io_cache_xcpt_pf_ld,
    input  io_cache_xcpt_pf_st,
    //output io_cache_invalidate_lr
    input  io_cache_ordered
);

  wire T0;
  wire T1;
  wire replaying_cmb;
  wire T2;
  wire T3;
  reg  replaying;
  wire T23;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg  R9;
  reg  R10;
  reg  s2_req_fire;
  reg  s1_req_fire;
  wire s0_req_fire;
  wire T11;
  wire T12;
  reg  s3_nack;
  wire[63:0] T13;
  wire[2:0] T14;
  wire[4:0] T15;
  wire[9:0] T16;
  wire[39:0] T17;
  wire T18;
  reg [63:0] R19;
  wire[63:0] T20;
  wire T21;
  wire T22;
  wire replayq1_io_deq_valid;
  wire[39:0] replayq1_io_deq_bits_addr;
  wire[9:0] replayq1_io_deq_bits_tag;
  wire[4:0] replayq1_io_deq_bits_cmd;
  wire[2:0] replayq1_io_deq_bits_typ;
  wire replayq1_io_deq_bits_kill;
  wire replayq1_io_deq_bits_phys;
  wire[63:0] replayq1_io_deq_bits_data;
  wire replayq2_io_deq_valid;
  wire[39:0] replayq2_io_deq_bits_addr;
  wire[9:0] replayq2_io_deq_bits_tag;
  wire[4:0] replayq2_io_deq_bits_cmd;
  wire[2:0] replayq2_io_deq_bits_typ;
  wire[63:0] replayq2_io_deq_bits_data;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire[39:0] req_arb_io_out_bits_addr;
  wire[9:0] req_arb_io_out_bits_tag;
  wire[4:0] req_arb_io_out_bits_cmd;
  wire[2:0] req_arb_io_out_bits_typ;
  wire[63:0] req_arb_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    replaying = {1{$random}};
    R9 = {1{$random}};
    R10 = {1{$random}};
    s2_req_fire = {1{$random}};
    s1_req_fire = {1{$random}};
    s3_nack = {1{$random}};
    R19 = {2{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_cache_invalidate_lr = {1{$random}};
//  assign io_requestor_ordered = {1{$random}};
//  assign io_requestor_xcpt_pf_st = {1{$random}};
//  assign io_requestor_xcpt_pf_ld = {1{$random}};
//  assign io_requestor_xcpt_ma_st = {1{$random}};
//  assign io_requestor_xcpt_ma_ld = {1{$random}};
//  assign io_requestor_replay_next_bits = {1{$random}};
//  assign io_requestor_replay_next_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T1 & io_requestor_req_valid;
  assign T1 = replaying_cmb ^ 1'h1;
  assign replaying_cmb = T2;
  assign T2 = T4 ? 1'h0 : T3;
  assign T3 = io_cache_resp_bits_nack ? 1'h1 : replaying;
  assign T23 = reset ? 1'h0 : replaying_cmb;
  assign T4 = T6 & T5;
  assign T5 = replayq2_io_deq_valid ^ 1'h1;
  assign T6 = T8 & T7;
  assign T7 = io_cache_resp_bits_nack ^ 1'h1;
  assign T8 = s2_req_fire & R9;
  assign s0_req_fire = io_cache_req_ready & io_cache_req_valid;
  assign T11 = T6 & replayq2_io_deq_valid;
  assign T12 = s2_req_fire & s3_nack;
  assign T13 = T11 ? replayq2_io_deq_bits_data : io_cache_resp_bits_store_data;
  assign T14 = T11 ? replayq2_io_deq_bits_typ : io_cache_resp_bits_typ;
  assign T15 = T11 ? replayq2_io_deq_bits_cmd : io_cache_resp_bits_cmd;
  assign T16 = T11 ? replayq2_io_deq_bits_tag : io_cache_resp_bits_tag;
  assign T17 = T11 ? replayq2_io_deq_bits_addr : io_cache_resp_bits_addr;
  assign T18 = T11 ? 1'h1 : io_cache_resp_bits_nack;
  assign io_cache_req_bits_data = R19;
  assign T20 = s0_req_fire ? req_arb_io_out_bits_data : R19;
  assign io_cache_req_bits_phys = 1'h1;
  assign io_cache_req_bits_kill = io_cache_resp_bits_nack;
  assign io_cache_req_bits_typ = req_arb_io_out_bits_typ;
  assign io_cache_req_bits_cmd = req_arb_io_out_bits_cmd;
  assign io_cache_req_bits_tag = req_arb_io_out_bits_tag;
  assign io_cache_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_cache_req_valid = req_arb_io_out_valid;
  assign io_requestor_resp_bits_store_data = io_cache_resp_bits_store_data;
  assign io_requestor_resp_bits_data_word_bypass = io_cache_resp_bits_data_word_bypass;
  assign io_requestor_resp_bits_has_data = io_cache_resp_bits_has_data;
  assign io_requestor_resp_bits_replay = io_cache_resp_bits_replay;
  assign io_requestor_resp_bits_nack = io_cache_resp_bits_nack;
  assign io_requestor_resp_bits_data = io_cache_resp_bits_data;
  assign io_requestor_resp_bits_typ = io_cache_resp_bits_typ;
  assign io_requestor_resp_bits_cmd = io_cache_resp_bits_cmd;
  assign io_requestor_resp_bits_tag = io_cache_resp_bits_tag;
  assign io_requestor_resp_bits_addr = io_cache_resp_bits_addr;
  assign io_requestor_resp_valid = io_cache_resp_valid;
  assign io_requestor_req_ready = T21;
  assign T21 = T22 & req_arb_io_in_1_ready;
  assign T22 = replaying_cmb ^ 1'h1;
  Queue_11 replayq1(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( T18 ),
       .io_enq_bits_addr( T17 ),
       .io_enq_bits_tag( T16 ),
       .io_enq_bits_cmd( T15 ),
       .io_enq_bits_typ( T14 ),
       //.io_enq_bits_kill(  )
       //.io_enq_bits_phys(  )
       .io_enq_bits_data( T13 ),
       .io_deq_ready( req_arb_io_in_0_ready ),
       .io_deq_valid( replayq1_io_deq_valid ),
       .io_deq_bits_addr( replayq1_io_deq_bits_addr ),
       .io_deq_bits_tag( replayq1_io_deq_bits_tag ),
       .io_deq_bits_cmd( replayq1_io_deq_bits_cmd ),
       .io_deq_bits_typ( replayq1_io_deq_bits_typ ),
       .io_deq_bits_kill( replayq1_io_deq_bits_kill ),
       .io_deq_bits_phys( replayq1_io_deq_bits_phys ),
       .io_deq_bits_data( replayq1_io_deq_bits_data )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign replayq1.io_enq_bits_kill = {1{$random}};
    assign replayq1.io_enq_bits_phys = {1{$random}};
// synthesis translate_on
`endif
  Queue_12 replayq2(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( T12 ),
       .io_enq_bits_addr( io_cache_resp_bits_addr ),
       .io_enq_bits_tag( io_cache_resp_bits_tag ),
       .io_enq_bits_cmd( io_cache_resp_bits_cmd ),
       .io_enq_bits_typ( io_cache_resp_bits_typ ),
       //.io_enq_bits_kill(  )
       //.io_enq_bits_phys(  )
       .io_enq_bits_data( io_cache_resp_bits_store_data ),
       .io_deq_ready( T11 ),
       .io_deq_valid( replayq2_io_deq_valid ),
       .io_deq_bits_addr( replayq2_io_deq_bits_addr ),
       .io_deq_bits_tag( replayq2_io_deq_bits_tag ),
       .io_deq_bits_cmd( replayq2_io_deq_bits_cmd ),
       .io_deq_bits_typ( replayq2_io_deq_bits_typ ),
       //.io_deq_bits_kill(  )
       //.io_deq_bits_phys(  )
       .io_deq_bits_data( replayq2_io_deq_bits_data )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign replayq2.io_enq_bits_kill = {1{$random}};
    assign replayq2.io_enq_bits_phys = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_5 req_arb(
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( T0 ),
       .io_in_1_bits_addr( io_requestor_req_bits_addr ),
       .io_in_1_bits_tag( io_requestor_req_bits_tag ),
       .io_in_1_bits_cmd( io_requestor_req_bits_cmd ),
       .io_in_1_bits_typ( io_requestor_req_bits_typ ),
       .io_in_1_bits_kill( io_requestor_req_bits_kill ),
       .io_in_1_bits_phys( io_requestor_req_bits_phys ),
       .io_in_1_bits_data( io_requestor_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( replayq1_io_deq_valid ),
       .io_in_0_bits_addr( replayq1_io_deq_bits_addr ),
       .io_in_0_bits_tag( replayq1_io_deq_bits_tag ),
       .io_in_0_bits_cmd( replayq1_io_deq_bits_cmd ),
       .io_in_0_bits_typ( replayq1_io_deq_bits_typ ),
       .io_in_0_bits_kill( replayq1_io_deq_bits_kill ),
       .io_in_0_bits_phys( replayq1_io_deq_bits_phys ),
       .io_in_0_bits_data( replayq1_io_deq_bits_data ),
       .io_out_ready( io_cache_req_ready ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_tag( req_arb_io_out_bits_tag ),
       .io_out_bits_cmd( req_arb_io_out_bits_cmd ),
       .io_out_bits_typ( req_arb_io_out_bits_typ ),
       //.io_out_bits_kill(  )
       //.io_out_bits_phys(  )
       .io_out_bits_data( req_arb_io_out_bits_data )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      replaying <= 1'h0;
    end else begin
      replaying <= replaying_cmb;
    end
    R9 <= R10;
    R10 <= replaying_cmb;
    s2_req_fire <= s1_req_fire;
    s1_req_fire <= s0_req_fire;
    s3_nack <= io_cache_resp_bits_nack;
    if(s0_req_fire) begin
      R19 <= req_arb_io_out_bits_data;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [4:0] io_enq_bits_rd,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[4:0] io_deq_bits_rd,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[68:0] T11;
  reg [68:0] ram [1:0];
  wire[68:0] T12;
  wire[68:0] T13;
  wire[68:0] T14;
  wire[4:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rd, io_enq_bits_data};
  assign io_deq_bits_rd = T15;
  assign T15 = T11[7'h44:7'h40];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module RocketTile(input clk, input reset,
    input  io_cached_0_acquire_ready,
    output io_cached_0_acquire_valid,
    output[25:0] io_cached_0_acquire_bits_addr_block,
    output[5:0] io_cached_0_acquire_bits_client_xact_id,
    output[1:0] io_cached_0_acquire_bits_addr_beat,
    output io_cached_0_acquire_bits_is_builtin_type,
    output[2:0] io_cached_0_acquire_bits_a_type,
    output[16:0] io_cached_0_acquire_bits_union,
    output[127:0] io_cached_0_acquire_bits_data,
    output io_cached_0_grant_ready,
    input  io_cached_0_grant_valid,
    input [1:0] io_cached_0_grant_bits_addr_beat,
    input [5:0] io_cached_0_grant_bits_client_xact_id,
    input [3:0] io_cached_0_grant_bits_manager_xact_id,
    input  io_cached_0_grant_bits_is_builtin_type,
    input [3:0] io_cached_0_grant_bits_g_type,
    input [127:0] io_cached_0_grant_bits_data,
    output io_cached_0_probe_ready,
    input  io_cached_0_probe_valid,
    input [25:0] io_cached_0_probe_bits_addr_block,
    input [1:0] io_cached_0_probe_bits_p_type,
    input  io_cached_0_release_ready,
    output io_cached_0_release_valid,
    output[1:0] io_cached_0_release_bits_addr_beat,
    output[25:0] io_cached_0_release_bits_addr_block,
    output[5:0] io_cached_0_release_bits_client_xact_id,
    output io_cached_0_release_bits_voluntary,
    output[2:0] io_cached_0_release_bits_r_type,
    output[127:0] io_cached_0_release_bits_data,
    input  io_uncached_0_acquire_ready,
    output io_uncached_0_acquire_valid,
    output[25:0] io_uncached_0_acquire_bits_addr_block,
    output[5:0] io_uncached_0_acquire_bits_client_xact_id,
    output[1:0] io_uncached_0_acquire_bits_addr_beat,
    output io_uncached_0_acquire_bits_is_builtin_type,
    output[2:0] io_uncached_0_acquire_bits_a_type,
    output[16:0] io_uncached_0_acquire_bits_union,
    output[127:0] io_uncached_0_acquire_bits_data,
    output io_uncached_0_grant_ready,
    input  io_uncached_0_grant_valid,
    input [1:0] io_uncached_0_grant_bits_addr_beat,
    input [5:0] io_uncached_0_grant_bits_client_xact_id,
    input [3:0] io_uncached_0_grant_bits_manager_xact_id,
    input  io_uncached_0_grant_bits_is_builtin_type,
    input [3:0] io_uncached_0_grant_bits_g_type,
    input [127:0] io_uncached_0_grant_bits_data,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    //input  io_dma_req_ready
    //output io_dma_req_valid
    //output[1:0] io_dma_req_bits_xact_id
    //output io_dma_req_bits_client_id
    //output[2:0] io_dma_req_bits_cmd
    //output[31:0] io_dma_req_bits_source
    //output[31:0] io_dma_req_bits_dest
    //output[31:0] io_dma_req_bits_length
    //output[1:0] io_dma_req_bits_size
    //output io_dma_resp_ready
    //input  io_dma_resp_valid
    //input [1:0] io_dma_resp_bits_xact_id
    //input  io_dma_resp_bits_client_id
    //input [1:0] io_dma_resp_bits_status
    input  init
);

  wire T0;
  wire dcArb_io_requestor_2_req_ready;
  wire dcArb_io_requestor_2_resp_valid;
  wire[39:0] dcArb_io_requestor_2_resp_bits_addr;
  wire[9:0] dcArb_io_requestor_2_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_2_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_2_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_2_resp_bits_data;
  wire dcArb_io_requestor_2_resp_bits_nack;
  wire dcArb_io_requestor_2_resp_bits_replay;
  wire dcArb_io_requestor_2_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_2_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_2_resp_bits_store_data;
  wire dcArb_io_requestor_2_replay_next_valid;
  wire[9:0] dcArb_io_requestor_2_replay_next_bits;
  wire dcArb_io_requestor_2_xcpt_ma_ld;
  wire dcArb_io_requestor_2_xcpt_ma_st;
  wire dcArb_io_requestor_2_xcpt_pf_ld;
  wire dcArb_io_requestor_2_xcpt_pf_st;
  wire dcArb_io_requestor_2_ordered;
  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[9:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[9:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[9:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[9:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire[39:0] dcArb_io_mem_req_bits_addr;
  wire[9:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_kill;
  wire dcArb_io_mem_req_bits_phys;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[4:0] RRArbiter_io_out_bits_rd;
  wire[63:0] RRArbiter_io_out_bits_data;
  wire SampleAccel_io_cmd_ready;
  wire SampleAccel_io_resp_valid;
  wire[4:0] SampleAccel_io_resp_bits_rd;
  wire[63:0] SampleAccel_io_resp_bits_data;
  wire SampleAccel_io_mem_req_valid;
  wire SampleAccel_io_mem_req_bits_phys;
  wire SampleAccel_io_busy;
  wire SampleAccel_io_interrupt;
  wire SampleAccel_io_autl_acquire_valid;
  wire SampleAccel_io_autl_grant_ready;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[4:0] Queue_io_deq_bits_rd;
  wire[63:0] Queue_io_deq_bits_data;
  wire core_io_host_csr_req_ready;
  wire core_io_host_csr_resp_valid;
  wire[63:0] core_io_host_csr_resp_bits;
  wire core_io_host_debug_stats_csr;
  wire core_io_imem_req_valid;
  wire[39:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_bits_mask;
  wire core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_btb_update_bits_pc;
  wire[38:0] core_io_imem_btb_update_bits_target;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isReturn;
  wire[38:0] core_io_imem_btb_update_bits_br_pc;
  wire core_io_imem_bht_update_valid;
  wire core_io_imem_bht_update_bits_prediction_valid;
  wire core_io_imem_bht_update_bits_prediction_bits_taken;
  wire core_io_imem_bht_update_bits_prediction_bits_mask;
  wire core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_bht_update_bits_pc;
  wire core_io_imem_bht_update_bits_taken;
  wire core_io_imem_bht_update_bits_mispredict;
  wire core_io_imem_ras_update_valid;
  wire core_io_imem_ras_update_bits_isCall;
  wire core_io_imem_ras_update_bits_isReturn;
  wire[38:0] core_io_imem_ras_update_bits_returnAddr;
  wire core_io_imem_ras_update_bits_prediction_valid;
  wire core_io_imem_ras_update_bits_prediction_bits_taken;
  wire core_io_imem_ras_update_bits_prediction_bits_mask;
  wire core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire[39:0] core_io_dmem_req_bits_addr;
  wire[9:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_bits_phys;
  wire[63:0] core_io_dmem_req_bits_data;
  wire core_io_dmem_invalidate_lr;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_status_sd;
  wire[30:0] core_io_ptw_status_zero2;
  wire core_io_ptw_status_sd_rv32;
  wire[8:0] core_io_ptw_status_zero1;
  wire[4:0] core_io_ptw_status_vm;
  wire core_io_ptw_status_mprv;
  wire[1:0] core_io_ptw_status_xs;
  wire[1:0] core_io_ptw_status_fs;
  wire[1:0] core_io_ptw_status_prv3;
  wire core_io_ptw_status_ie3;
  wire[1:0] core_io_ptw_status_prv2;
  wire core_io_ptw_status_ie2;
  wire[1:0] core_io_ptw_status_prv1;
  wire core_io_ptw_status_ie1;
  wire[1:0] core_io_ptw_status_prv;
  wire core_io_ptw_status_ie;
  wire[31:0] core_io_fpu_inst;
  wire[63:0] core_io_fpu_fromint_data;
  wire[2:0] core_io_fpu_fcsr_rm;
  wire core_io_fpu_dmem_resp_val;
  wire[2:0] core_io_fpu_dmem_resp_type;
  wire[4:0] core_io_fpu_dmem_resp_tag;
  wire[63:0] core_io_fpu_dmem_resp_data;
  wire core_io_fpu_valid;
  wire core_io_fpu_killx;
  wire core_io_fpu_killm;
  wire core_io_rocc_cmd_valid;
  wire[6:0] core_io_rocc_cmd_bits_inst_funct;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire core_io_rocc_cmd_bits_inst_xd;
  wire core_io_rocc_cmd_bits_inst_xs1;
  wire core_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] core_io_rocc_cmd_bits_inst_rd;
  wire[6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] core_io_rocc_cmd_bits_rs1;
  wire[63:0] core_io_rocc_cmd_bits_rs2;
  wire core_io_rocc_resp_ready;
  wire core_io_rocc_s;
  wire core_io_rocc_exception;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[19:0] ptw_io_requestor_1_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_1_resp_bits_pte_d;
  wire ptw_io_requestor_1_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_1_resp_bits_pte_typ;
  wire ptw_io_requestor_1_resp_bits_pte_v;
  wire ptw_io_requestor_1_status_sd;
  wire[30:0] ptw_io_requestor_1_status_zero2;
  wire ptw_io_requestor_1_status_sd_rv32;
  wire[8:0] ptw_io_requestor_1_status_zero1;
  wire[4:0] ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_mprv;
  wire[1:0] ptw_io_requestor_1_status_xs;
  wire[1:0] ptw_io_requestor_1_status_fs;
  wire[1:0] ptw_io_requestor_1_status_prv3;
  wire ptw_io_requestor_1_status_ie3;
  wire[1:0] ptw_io_requestor_1_status_prv2;
  wire ptw_io_requestor_1_status_ie2;
  wire[1:0] ptw_io_requestor_1_status_prv1;
  wire ptw_io_requestor_1_status_ie1;
  wire[1:0] ptw_io_requestor_1_status_prv;
  wire ptw_io_requestor_1_status_ie;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[19:0] ptw_io_requestor_0_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_0_resp_bits_pte_d;
  wire ptw_io_requestor_0_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_0_resp_bits_pte_typ;
  wire ptw_io_requestor_0_resp_bits_pte_v;
  wire ptw_io_requestor_0_status_sd;
  wire[30:0] ptw_io_requestor_0_status_zero2;
  wire ptw_io_requestor_0_status_sd_rv32;
  wire[8:0] ptw_io_requestor_0_status_zero1;
  wire[4:0] ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_mprv;
  wire[1:0] ptw_io_requestor_0_status_xs;
  wire[1:0] ptw_io_requestor_0_status_fs;
  wire[1:0] ptw_io_requestor_0_status_prv3;
  wire ptw_io_requestor_0_status_ie3;
  wire[1:0] ptw_io_requestor_0_status_prv2;
  wire ptw_io_requestor_0_status_ie2;
  wire[1:0] ptw_io_requestor_0_status_prv1;
  wire ptw_io_requestor_0_status_ie1;
  wire[1:0] ptw_io_requestor_0_status_prv;
  wire ptw_io_requestor_0_status_ie;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_mem_req_valid;
  wire[39:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_bits_phys;
  wire[63:0] ptw_io_mem_req_bits_data;
  wire ClientTileLinkIOArbiter_io_in_1_acquire_ready;
  wire ClientTileLinkIOArbiter_io_in_1_grant_valid;
  wire[1:0] ClientTileLinkIOArbiter_io_in_1_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkIOArbiter_io_in_1_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOArbiter_io_in_1_grant_bits_manager_xact_id;
  wire ClientTileLinkIOArbiter_io_in_1_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOArbiter_io_in_1_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOArbiter_io_in_1_grant_bits_data;
  wire ClientTileLinkIOArbiter_io_in_0_acquire_ready;
  wire ClientTileLinkIOArbiter_io_in_0_grant_valid;
  wire[1:0] ClientTileLinkIOArbiter_io_in_0_grant_bits_addr_beat;
  wire[5:0] ClientTileLinkIOArbiter_io_in_0_grant_bits_client_xact_id;
  wire[3:0] ClientTileLinkIOArbiter_io_in_0_grant_bits_manager_xact_id;
  wire ClientTileLinkIOArbiter_io_in_0_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOArbiter_io_in_0_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOArbiter_io_in_0_grant_bits_data;
  wire ClientTileLinkIOArbiter_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOArbiter_io_out_acquire_bits_addr_block;
  wire[5:0] ClientTileLinkIOArbiter_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOArbiter_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOArbiter_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOArbiter_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOArbiter_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOArbiter_io_out_acquire_bits_data;
  wire ClientTileLinkIOArbiter_io_out_grant_ready;
  wire RoccCommandRouter_io_in_ready;
  wire RoccCommandRouter_io_out_0_valid;
  wire[6:0] RoccCommandRouter_io_out_0_bits_inst_funct;
  wire[4:0] RoccCommandRouter_io_out_0_bits_inst_rs2;
  wire[4:0] RoccCommandRouter_io_out_0_bits_inst_rs1;
  wire RoccCommandRouter_io_out_0_bits_inst_xd;
  wire RoccCommandRouter_io_out_0_bits_inst_xs1;
  wire RoccCommandRouter_io_out_0_bits_inst_xs2;
  wire[4:0] RoccCommandRouter_io_out_0_bits_inst_rd;
  wire[6:0] RoccCommandRouter_io_out_0_bits_inst_opcode;
  wire[63:0] RoccCommandRouter_io_out_0_bits_rs1;
  wire[63:0] RoccCommandRouter_io_out_0_bits_rs2;
  wire RoccCommandRouter_io_busy;
  wire SimpleHellaCacheIF_io_requestor_req_ready;
  wire SimpleHellaCacheIF_io_requestor_resp_valid;
  
  wire [39:0] SimpleHellaCacheIF_io_requestor_req_addr;
  wire [9:0] SimpleHellaCacheIF_io_requestor_req_tag;
  wire [4:0] SimpleHellaCacheIF_io_requestor_req_cmd;
  wire [2:0] SimpleHellaCacheIF_io_requestor_req_typ;
  wire SimpleHellaCacheIF_io_requestor_req_kill;
  wire SimpleHellaCacheIF_io_requestor_req_phys;
  wire [63:0] SimpleHellaCacheIF_io_requestor_req_data;
  
  wire[39:0] SimpleHellaCacheIF_io_requestor_resp_bits_addr;
  wire[9:0] SimpleHellaCacheIF_io_requestor_resp_bits_tag;
  wire[4:0] SimpleHellaCacheIF_io_requestor_resp_bits_cmd;
  wire[2:0] SimpleHellaCacheIF_io_requestor_resp_bits_typ;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_data;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_nack;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_replay;
  wire SimpleHellaCacheIF_io_requestor_resp_bits_has_data;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_data_word_bypass;
  wire[63:0] SimpleHellaCacheIF_io_requestor_resp_bits_store_data;
  wire SimpleHellaCacheIF_io_cache_req_valid;
  wire[39:0] SimpleHellaCacheIF_io_cache_req_bits_addr;
  wire[9:0] SimpleHellaCacheIF_io_cache_req_bits_tag;
  wire[4:0] SimpleHellaCacheIF_io_cache_req_bits_cmd;
  wire[2:0] SimpleHellaCacheIF_io_cache_req_bits_typ;
  wire SimpleHellaCacheIF_io_cache_req_bits_kill;
  wire SimpleHellaCacheIF_io_cache_req_bits_phys;
  wire[63:0] SimpleHellaCacheIF_io_cache_req_bits_data;
  wire icache_io_cpu_resp_valid;
  wire[39:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data_0;
  wire icache_io_cpu_resp_bits_mask;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_bits_mask;
  wire icache_io_cpu_btb_resp_bits_bridx;
  wire[38:0] icache_io_cpu_btb_resp_bits_target;
  wire[5:0] icache_io_cpu_btb_resp_bits_entry;
  wire[6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[39:0] icache_io_cpu_npc;
  wire icache_io_ptw_req_valid;
  wire[26:0] icache_io_ptw_req_bits_addr;
  wire[1:0] icache_io_ptw_req_bits_prv;
  wire icache_io_ptw_req_bits_store;
  wire icache_io_ptw_req_bits_fetch;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[5:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[39:0] dcache_io_cpu_resp_bits_addr;
  wire[9:0] dcache_io_cpu_resp_bits_tag;
  wire[4:0] dcache_io_cpu_resp_bits_cmd;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_word_bypass;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[9:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ordered;
  wire dcache_io_ptw_req_valid;
  wire[26:0] dcache_io_ptw_req_bits_addr;
  wire[1:0] dcache_io_ptw_req_bits_prv;
  wire dcache_io_ptw_req_bits_store;
  wire dcache_io_ptw_req_bits_fetch;
  wire dcache_io_mem_acquire_valid;
  wire[25:0] dcache_io_mem_acquire_bits_addr_block;
  wire[5:0] dcache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] dcache_io_mem_acquire_bits_addr_beat;
  wire dcache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] dcache_io_mem_acquire_bits_a_type;
  wire[16:0] dcache_io_mem_acquire_bits_union;
  wire[127:0] dcache_io_mem_acquire_bits_data;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_addr_beat;
  wire[25:0] dcache_io_mem_release_bits_addr_block;
  wire[5:0] dcache_io_mem_release_bits_client_xact_id;
  wire dcache_io_mem_release_bits_voluntary;
  wire[2:0] dcache_io_mem_release_bits_r_type;
  wire[127:0] dcache_io_mem_release_bits_data;
  wire FPU_io_fcsr_flags_valid;
  wire[4:0] FPU_io_fcsr_flags_bits;
  wire[63:0] FPU_io_store_data;
  wire[63:0] FPU_io_toint_data;
  wire FPU_io_fcsr_rdy;
  wire FPU_io_nack_mem;
  wire FPU_io_illegal_rm;
  wire[4:0] FPU_io_dec_cmd;
  wire FPU_io_dec_ldst;
  wire FPU_io_dec_wen;
  wire FPU_io_dec_ren1;
  wire FPU_io_dec_ren2;
  wire FPU_io_dec_ren3;
  wire FPU_io_dec_swap12;
  wire FPU_io_dec_swap23;
  wire FPU_io_dec_single;
  wire FPU_io_dec_fromint;
  wire FPU_io_dec_toint;
  wire FPU_io_dec_fastpipe;
  wire FPU_io_dec_fma;
  wire FPU_io_dec_div;
  wire FPU_io_dec_sqrt;
  wire FPU_io_dec_round;
  wire FPU_io_dec_wflags;
  wire FPU_io_sboard_set;
  wire FPU_io_sboard_clr;
  wire[4:0] FPU_io_sboard_clra;
  wire FPU_io_cp_req_ready;
  wire FPU_io_cp_resp_valid;
  wire[64:0] FPU_io_cp_resp_bits_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_dma_resp_ready = {1{$random}};
//  assign io_dma_req_bits_size = {1{$random}};
//  assign io_dma_req_bits_length = {1{$random}};
//  assign io_dma_req_bits_dest = {1{$random}};
//  assign io_dma_req_bits_source = {1{$random}};
//  assign io_dma_req_bits_cmd = {1{$random}};
//  assign io_dma_req_bits_client_id = {1{$random}};
//  assign io_dma_req_bits_xact_id = {1{$random}};
//  assign io_dma_req_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = RoccCommandRouter_io_busy | SampleAccel_io_busy;
  assign io_host_debug_stats_csr = core_io_host_debug_stats_csr;
  assign io_host_csr_resp_bits = core_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = core_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = core_io_host_csr_req_ready;
  assign io_uncached_0_grant_ready = ClientTileLinkIOArbiter_io_out_grant_ready;
  assign io_uncached_0_acquire_bits_data = ClientTileLinkIOArbiter_io_out_acquire_bits_data;
  assign io_uncached_0_acquire_bits_union = ClientTileLinkIOArbiter_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_a_type = ClientTileLinkIOArbiter_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_is_builtin_type = ClientTileLinkIOArbiter_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_addr_beat = ClientTileLinkIOArbiter_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_client_xact_id = ClientTileLinkIOArbiter_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_block = ClientTileLinkIOArbiter_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_valid = ClientTileLinkIOArbiter_io_out_acquire_valid;
  assign io_cached_0_release_bits_data = dcache_io_mem_release_bits_data;
  assign io_cached_0_release_bits_r_type = dcache_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_voluntary = dcache_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_client_xact_id = dcache_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_addr_block = dcache_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_addr_beat = dcache_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_valid = dcache_io_mem_release_valid;
  assign io_cached_0_probe_ready = dcache_io_mem_probe_ready;
  assign io_cached_0_grant_ready = dcache_io_mem_grant_ready;
  assign io_cached_0_acquire_bits_data = dcache_io_mem_acquire_bits_data;
  assign io_cached_0_acquire_bits_union = dcache_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_a_type = dcache_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_is_builtin_type = dcache_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_addr_beat = dcache_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_client_xact_id = dcache_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_block = dcache_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_valid = dcache_io_mem_acquire_valid;
  Rocket core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( core_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( core_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( core_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( core_io_host_debug_stats_csr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_imem_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_imem_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_imem_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_imem_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_imem_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_imem_npc( icache_io_cpu_npc ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_dmem_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_status_sd( core_io_ptw_status_sd ),
       .io_ptw_status_zero2( core_io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( core_io_ptw_status_zero1 ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_mprv( core_io_ptw_status_mprv ),
       .io_ptw_status_xs( core_io_ptw_status_xs ),
       .io_ptw_status_fs( core_io_ptw_status_fs ),
       .io_ptw_status_prv3( core_io_ptw_status_prv3 ),
       .io_ptw_status_ie3( core_io_ptw_status_ie3 ),
       .io_ptw_status_prv2( core_io_ptw_status_prv2 ),
       .io_ptw_status_ie2( core_io_ptw_status_ie2 ),
       .io_ptw_status_prv1( core_io_ptw_status_prv1 ),
       .io_ptw_status_ie1( core_io_ptw_status_ie1 ),
       .io_ptw_status_prv( core_io_ptw_status_prv ),
       .io_ptw_status_ie( core_io_ptw_status_ie ),
       .io_fpu_inst( core_io_fpu_inst ),
       .io_fpu_fromint_data( core_io_fpu_fromint_data ),
       .io_fpu_fcsr_rm( core_io_fpu_fcsr_rm ),
       .io_fpu_fcsr_flags_valid( FPU_io_fcsr_flags_valid ),
       .io_fpu_fcsr_flags_bits( FPU_io_fcsr_flags_bits ),
       .io_fpu_store_data( FPU_io_store_data ),
       .io_fpu_toint_data( FPU_io_toint_data ),
       .io_fpu_dmem_resp_val( core_io_fpu_dmem_resp_val ),
       .io_fpu_dmem_resp_type( core_io_fpu_dmem_resp_type ),
       .io_fpu_dmem_resp_tag( core_io_fpu_dmem_resp_tag ),
       .io_fpu_dmem_resp_data( core_io_fpu_dmem_resp_data ),
       .io_fpu_valid( core_io_fpu_valid ),
       .io_fpu_fcsr_rdy( FPU_io_fcsr_rdy ),
       .io_fpu_nack_mem( FPU_io_nack_mem ),
       .io_fpu_illegal_rm( FPU_io_illegal_rm ),
       .io_fpu_killx( core_io_fpu_killx ),
       .io_fpu_killm( core_io_fpu_killm ),
       .io_fpu_dec_cmd( FPU_io_dec_cmd ),
       .io_fpu_dec_ldst( FPU_io_dec_ldst ),
       .io_fpu_dec_wen( FPU_io_dec_wen ),
       .io_fpu_dec_ren1( FPU_io_dec_ren1 ),
       .io_fpu_dec_ren2( FPU_io_dec_ren2 ),
       .io_fpu_dec_ren3( FPU_io_dec_ren3 ),
       .io_fpu_dec_swap12( FPU_io_dec_swap12 ),
       .io_fpu_dec_swap23( FPU_io_dec_swap23 ),
       .io_fpu_dec_single( FPU_io_dec_single ),
       .io_fpu_dec_fromint( FPU_io_dec_fromint ),
       .io_fpu_dec_toint( FPU_io_dec_toint ),
       .io_fpu_dec_fastpipe( FPU_io_dec_fastpipe ),
       .io_fpu_dec_fma( FPU_io_dec_fma ),
       .io_fpu_dec_div( FPU_io_dec_div ),
       .io_fpu_dec_sqrt( FPU_io_dec_sqrt ),
       .io_fpu_dec_round( FPU_io_dec_round ),
       .io_fpu_dec_wflags( FPU_io_dec_wflags ),
       .io_fpu_sboard_set( FPU_io_sboard_set ),
       .io_fpu_sboard_clr( FPU_io_sboard_clr ),
       .io_fpu_sboard_clra( FPU_io_sboard_clra ),
       .io_fpu_cp_req_ready( FPU_io_cp_req_ready ),
       //.io_fpu_cp_req_valid(  )
       //.io_fpu_cp_req_bits_cmd(  )
       //.io_fpu_cp_req_bits_ldst(  )
       //.io_fpu_cp_req_bits_wen(  )
       //.io_fpu_cp_req_bits_ren1(  )
       //.io_fpu_cp_req_bits_ren2(  )
       //.io_fpu_cp_req_bits_ren3(  )
       //.io_fpu_cp_req_bits_swap12(  )
       //.io_fpu_cp_req_bits_swap23(  )
       //.io_fpu_cp_req_bits_single(  )
       //.io_fpu_cp_req_bits_fromint(  )
       //.io_fpu_cp_req_bits_toint(  )
       //.io_fpu_cp_req_bits_fastpipe(  )
       //.io_fpu_cp_req_bits_fma(  )
       //.io_fpu_cp_req_bits_div(  )
       //.io_fpu_cp_req_bits_sqrt(  )
       //.io_fpu_cp_req_bits_round(  )
       //.io_fpu_cp_req_bits_wflags(  )
       //.io_fpu_cp_req_bits_rm(  )
       //.io_fpu_cp_req_bits_typ(  )
       //.io_fpu_cp_req_bits_in1(  )
       //.io_fpu_cp_req_bits_in2(  )
       //.io_fpu_cp_req_bits_in3(  )
       //.io_fpu_cp_resp_ready(  )
       .io_fpu_cp_resp_valid( FPU_io_cp_resp_valid ),
       .io_fpu_cp_resp_bits_data( FPU_io_cp_resp_bits_data ),
       //.io_fpu_cp_resp_bits_exc(  )
       .io_rocc_cmd_ready( RoccCommandRouter_io_in_ready ),
       .io_rocc_cmd_valid( core_io_rocc_cmd_valid ),
       .io_rocc_cmd_bits_inst_funct( core_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( core_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( core_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( core_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( core_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( core_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( core_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( core_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( core_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( core_io_rocc_cmd_bits_rs2 ),
       .io_rocc_resp_ready( core_io_rocc_resp_ready ),
       .io_rocc_resp_valid( RRArbiter_io_out_valid ),
       .io_rocc_resp_bits_rd( RRArbiter_io_out_bits_rd ),
       .io_rocc_resp_bits_data( RRArbiter_io_out_bits_data ),
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_invalidate_lr(  )
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( T0 ),
       .io_rocc_s( core_io_rocc_s ),
       .io_rocc_interrupt( SampleAccel_io_interrupt ),
       //.io_rocc_autl_acquire_ready(  )
       //.io_rocc_autl_acquire_valid(  )
       //.io_rocc_autl_acquire_bits_addr_block(  )
       //.io_rocc_autl_acquire_bits_client_xact_id(  )
       //.io_rocc_autl_acquire_bits_addr_beat(  )
       //.io_rocc_autl_acquire_bits_is_builtin_type(  )
       //.io_rocc_autl_acquire_bits_a_type(  )
       //.io_rocc_autl_acquire_bits_union(  )
       //.io_rocc_autl_acquire_bits_data(  )
       //.io_rocc_autl_grant_ready(  )
       //.io_rocc_autl_grant_valid(  )
       //.io_rocc_autl_grant_bits_addr_beat(  )
       //.io_rocc_autl_grant_bits_client_xact_id(  )
       //.io_rocc_autl_grant_bits_manager_xact_id(  )
       //.io_rocc_autl_grant_bits_is_builtin_type(  )
       //.io_rocc_autl_grant_bits_g_type(  )
       //.io_rocc_autl_grant_bits_data(  )
       //.io_rocc_fpu_req_ready(  )
       //.io_rocc_fpu_req_valid(  )
       //.io_rocc_fpu_req_bits_cmd(  )
       //.io_rocc_fpu_req_bits_ldst(  )
       //.io_rocc_fpu_req_bits_wen(  )
       //.io_rocc_fpu_req_bits_ren1(  )
       //.io_rocc_fpu_req_bits_ren2(  )
       //.io_rocc_fpu_req_bits_ren3(  )
       //.io_rocc_fpu_req_bits_swap12(  )
       //.io_rocc_fpu_req_bits_swap23(  )
       //.io_rocc_fpu_req_bits_single(  )
       //.io_rocc_fpu_req_bits_fromint(  )
       //.io_rocc_fpu_req_bits_toint(  )
       //.io_rocc_fpu_req_bits_fastpipe(  )
       //.io_rocc_fpu_req_bits_fma(  )
       //.io_rocc_fpu_req_bits_div(  )
       //.io_rocc_fpu_req_bits_sqrt(  )
       //.io_rocc_fpu_req_bits_round(  )
       //.io_rocc_fpu_req_bits_wflags(  )
       //.io_rocc_fpu_req_bits_rm(  )
       //.io_rocc_fpu_req_bits_typ(  )
       //.io_rocc_fpu_req_bits_in1(  )
       //.io_rocc_fpu_req_bits_in2(  )
       //.io_rocc_fpu_req_bits_in3(  )
       //.io_rocc_fpu_resp_ready(  )
       //.io_rocc_fpu_resp_valid(  )
       //.io_rocc_fpu_resp_bits_data(  )
       //.io_rocc_fpu_resp_bits_exc(  )
       .io_rocc_exception( core_io_rocc_exception )
       //.io_rocc_csr_waddr(  )
       //.io_rocc_csr_wdata(  )
       //.io_rocc_csr_wen(  )
       //.io_rocc_host_id(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_invalidate_lr = {1{$random}};
    assign core.io_rocc_autl_acquire_valid = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_union = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_data = {4{$random}};
    assign core.io_rocc_autl_grant_ready = {1{$random}};
    assign core.io_rocc_fpu_req_valid = {1{$random}};
    assign core.io_rocc_fpu_req_bits_cmd = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ldst = {1{$random}};
    assign core.io_rocc_fpu_req_bits_wen = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren1 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren2 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren3 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_swap12 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_swap23 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_single = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fromint = {1{$random}};
    assign core.io_rocc_fpu_req_bits_toint = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fastpipe = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fma = {1{$random}};
    assign core.io_rocc_fpu_req_bits_div = {1{$random}};
    assign core.io_rocc_fpu_req_bits_sqrt = {1{$random}};
    assign core.io_rocc_fpu_req_bits_round = {1{$random}};
    assign core.io_rocc_fpu_req_bits_wflags = {1{$random}};
    assign core.io_rocc_fpu_req_bits_rm = {1{$random}};
    assign core.io_rocc_fpu_req_bits_typ = {1{$random}};
    assign core.io_rocc_fpu_req_bits_in1 = {3{$random}};
    assign core.io_rocc_fpu_req_bits_in2 = {3{$random}};
    assign core.io_rocc_fpu_req_bits_in3 = {3{$random}};
    assign core.io_rocc_fpu_resp_ready = {1{$random}};
// synthesis translate_on
`endif
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_cpu_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_cpu_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_cpu_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_cpu_btb_update_bits_taken(  )
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_cpu_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_cpu_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_cpu_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_cpu_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_cpu_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_cpu_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_cpu_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_cpu_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_cpu_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_cpu_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_cpu_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_cpu_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_cpu_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_cpu_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_cpu_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_cpu_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_cpu_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_cpu_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_cpu_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_cpu_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_cpu_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_cpu_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_cpu_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_cpu_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_cpu_npc( icache_io_cpu_npc ),
       .io_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_ptw_req_valid( icache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_0_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_0_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_0_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_0_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_0_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_acquire_ready( ClientTileLinkIOArbiter_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( ClientTileLinkIOArbiter_io_in_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( ClientTileLinkIOArbiter_io_in_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( ClientTileLinkIOArbiter_io_in_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( ClientTileLinkIOArbiter_io_in_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( ClientTileLinkIOArbiter_io_in_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( ClientTileLinkIOArbiter_io_in_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( ClientTileLinkIOArbiter_io_in_0_grant_bits_data ),
       .init( init )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign icache.io_cpu_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_ptw_req_valid( dcache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_1_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_1_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_1_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_1_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_1_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_mem_acquire_ready( io_cached_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( dcache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( dcache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( dcache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( dcache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( dcache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( dcache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( dcache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_cached_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_cached_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_cached_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_cached_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_cached_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_cached_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_cached_0_grant_bits_data ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_cached_0_probe_valid ),
       .io_mem_probe_bits_addr_block( io_cached_0_probe_bits_addr_block ),
       .io_mem_probe_bits_p_type( io_cached_0_probe_bits_p_type ),
       .io_mem_release_ready( io_cached_0_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_addr_beat( dcache_io_mem_release_bits_addr_beat ),
       .io_mem_release_bits_addr_block( dcache_io_mem_release_bits_addr_block ),
       .io_mem_release_bits_client_xact_id( dcache_io_mem_release_bits_client_xact_id ),
       .io_mem_release_bits_voluntary( dcache_io_mem_release_bits_voluntary ),
       .io_mem_release_bits_r_type( dcache_io_mem_release_bits_r_type ),
       .io_mem_release_bits_data( dcache_io_mem_release_bits_data ),
       .init( init )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_ptw_req_valid ),
       .io_requestor_1_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_requestor_1_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_requestor_1_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_requestor_1_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_requestor_1_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_requestor_1_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_requestor_1_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_requestor_1_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_requestor_1_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_requestor_1_status_sd( ptw_io_requestor_1_status_sd ),
       .io_requestor_1_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_requestor_1_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_requestor_1_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_requestor_1_status_xs( ptw_io_requestor_1_status_xs ),
       .io_requestor_1_status_fs( ptw_io_requestor_1_status_fs ),
       .io_requestor_1_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_requestor_1_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_requestor_1_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_requestor_1_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_requestor_1_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_requestor_1_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_requestor_1_status_prv( ptw_io_requestor_1_status_prv ),
       .io_requestor_1_status_ie( ptw_io_requestor_1_status_ie ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_ptw_req_valid ),
       .io_requestor_0_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_requestor_0_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_requestor_0_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_requestor_0_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_requestor_0_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_requestor_0_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_requestor_0_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_requestor_0_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_requestor_0_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_requestor_0_status_sd( ptw_io_requestor_0_status_sd ),
       .io_requestor_0_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_requestor_0_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_requestor_0_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_requestor_0_status_xs( ptw_io_requestor_0_status_xs ),
       .io_requestor_0_status_fs( ptw_io_requestor_0_status_fs ),
       .io_requestor_0_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_requestor_0_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_requestor_0_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_requestor_0_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_requestor_0_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_requestor_0_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_requestor_0_status_prv( ptw_io_requestor_0_status_prv ),
       .io_requestor_0_status_ie( ptw_io_requestor_0_status_ie ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_status_sd( core_io_ptw_status_sd ),
       .io_dpath_status_zero2( core_io_ptw_status_zero2 ),
       .io_dpath_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_dpath_status_zero1( core_io_ptw_status_zero1 ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_mprv( core_io_ptw_status_mprv ),
       .io_dpath_status_xs( core_io_ptw_status_xs ),
       .io_dpath_status_fs( core_io_ptw_status_fs ),
       .io_dpath_status_prv3( core_io_ptw_status_prv3 ),
       .io_dpath_status_ie3( core_io_ptw_status_ie3 ),
       .io_dpath_status_prv2( core_io_ptw_status_prv2 ),
       .io_dpath_status_ie2( core_io_ptw_status_ie2 ),
       .io_dpath_status_prv1( core_io_ptw_status_prv1 ),
       .io_dpath_status_ie1( core_io_ptw_status_ie1 ),
       .io_dpath_status_prv( core_io_ptw_status_prv ),
       .io_dpath_status_ie( core_io_ptw_status_ie )
  );
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_2_req_ready( dcArb_io_requestor_2_req_ready ),
       .io_requestor_2_req_valid( SimpleHellaCacheIF_io_cache_req_valid ),
       .io_requestor_2_req_bits_addr( SimpleHellaCacheIF_io_cache_req_bits_addr ),
       .io_requestor_2_req_bits_tag( SimpleHellaCacheIF_io_cache_req_bits_tag ),
       .io_requestor_2_req_bits_cmd( SimpleHellaCacheIF_io_cache_req_bits_cmd ),
       .io_requestor_2_req_bits_typ( SimpleHellaCacheIF_io_cache_req_bits_typ ),
       .io_requestor_2_req_bits_kill( SimpleHellaCacheIF_io_cache_req_bits_kill ),
       .io_requestor_2_req_bits_phys( SimpleHellaCacheIF_io_cache_req_bits_phys ),
       .io_requestor_2_req_bits_data( SimpleHellaCacheIF_io_cache_req_bits_data ),
       .io_requestor_2_resp_valid( dcArb_io_requestor_2_resp_valid ),
       .io_requestor_2_resp_bits_addr( dcArb_io_requestor_2_resp_bits_addr ),
       .io_requestor_2_resp_bits_tag( dcArb_io_requestor_2_resp_bits_tag ),
       .io_requestor_2_resp_bits_cmd( dcArb_io_requestor_2_resp_bits_cmd ),
       .io_requestor_2_resp_bits_typ( dcArb_io_requestor_2_resp_bits_typ ),
       .io_requestor_2_resp_bits_data( dcArb_io_requestor_2_resp_bits_data ),
       .io_requestor_2_resp_bits_nack( dcArb_io_requestor_2_resp_bits_nack ),
       .io_requestor_2_resp_bits_replay( dcArb_io_requestor_2_resp_bits_replay ),
       .io_requestor_2_resp_bits_has_data( dcArb_io_requestor_2_resp_bits_has_data ),
       .io_requestor_2_resp_bits_data_word_bypass( dcArb_io_requestor_2_resp_bits_data_word_bypass ),
       .io_requestor_2_resp_bits_store_data( dcArb_io_requestor_2_resp_bits_store_data ),
       .io_requestor_2_replay_next_valid( dcArb_io_requestor_2_replay_next_valid ),
       .io_requestor_2_replay_next_bits( dcArb_io_requestor_2_replay_next_bits ),
       .io_requestor_2_xcpt_ma_ld( dcArb_io_requestor_2_xcpt_ma_ld ),
       .io_requestor_2_xcpt_ma_st( dcArb_io_requestor_2_xcpt_ma_st ),
       .io_requestor_2_xcpt_pf_ld( dcArb_io_requestor_2_xcpt_pf_ld ),
       .io_requestor_2_xcpt_pf_st( dcArb_io_requestor_2_xcpt_pf_st ),
       //.io_requestor_2_invalidate_lr(  )
       .io_requestor_2_ordered( dcArb_io_requestor_2_ordered ),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_requestor_1_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_invalidate_lr(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
  FPU FPU(.clk(clk), .reset(reset),
       .io_inst( core_io_fpu_inst ),
       .io_fromint_data( core_io_fpu_fromint_data ),
       .io_fcsr_rm( core_io_fpu_fcsr_rm ),
       .io_fcsr_flags_valid( FPU_io_fcsr_flags_valid ),
       .io_fcsr_flags_bits( FPU_io_fcsr_flags_bits ),
       .io_store_data( FPU_io_store_data ),
       .io_toint_data( FPU_io_toint_data ),
       .io_dmem_resp_val( core_io_fpu_dmem_resp_val ),
       .io_dmem_resp_type( core_io_fpu_dmem_resp_type ),
       .io_dmem_resp_tag( core_io_fpu_dmem_resp_tag ),
       .io_dmem_resp_data( core_io_fpu_dmem_resp_data ),
       .io_valid( core_io_fpu_valid ),
       .io_fcsr_rdy( FPU_io_fcsr_rdy ),
       .io_nack_mem( FPU_io_nack_mem ),
       .io_illegal_rm( FPU_io_illegal_rm ),
       .io_killx( core_io_fpu_killx ),
       .io_killm( core_io_fpu_killm ),
       .io_dec_cmd( FPU_io_dec_cmd ),
       .io_dec_ldst( FPU_io_dec_ldst ),
       .io_dec_wen( FPU_io_dec_wen ),
       .io_dec_ren1( FPU_io_dec_ren1 ),
       .io_dec_ren2( FPU_io_dec_ren2 ),
       .io_dec_ren3( FPU_io_dec_ren3 ),
       .io_dec_swap12( FPU_io_dec_swap12 ),
       .io_dec_swap23( FPU_io_dec_swap23 ),
       .io_dec_single( FPU_io_dec_single ),
       .io_dec_fromint( FPU_io_dec_fromint ),
       .io_dec_toint( FPU_io_dec_toint ),
       .io_dec_fastpipe( FPU_io_dec_fastpipe ),
       .io_dec_fma( FPU_io_dec_fma ),
       .io_dec_div( FPU_io_dec_div ),
       .io_dec_sqrt( FPU_io_dec_sqrt ),
       .io_dec_round( FPU_io_dec_round ),
       .io_dec_wflags( FPU_io_dec_wflags ),
       .io_sboard_set( FPU_io_sboard_set ),
       .io_sboard_clr( FPU_io_sboard_clr ),
       .io_sboard_clra( FPU_io_sboard_clra ),
       .io_cp_req_ready( FPU_io_cp_req_ready ),
       .io_cp_req_valid( 1'h0 ),
       //.io_cp_req_bits_cmd(  )
       //.io_cp_req_bits_ldst(  )
       //.io_cp_req_bits_wen(  )
       //.io_cp_req_bits_ren1(  )
       //.io_cp_req_bits_ren2(  )
       //.io_cp_req_bits_ren3(  )
       //.io_cp_req_bits_swap12(  )
       //.io_cp_req_bits_swap23(  )
       //.io_cp_req_bits_single(  )
       //.io_cp_req_bits_fromint(  )
       //.io_cp_req_bits_toint(  )
       //.io_cp_req_bits_fastpipe(  )
       //.io_cp_req_bits_fma(  )
       //.io_cp_req_bits_div(  )
       //.io_cp_req_bits_sqrt(  )
       //.io_cp_req_bits_round(  )
       //.io_cp_req_bits_wflags(  )
       //.io_cp_req_bits_rm(  )
       //.io_cp_req_bits_typ(  )
       //.io_cp_req_bits_in1(  )
       //.io_cp_req_bits_in2(  )
       //.io_cp_req_bits_in3(  )
       .io_cp_resp_ready( 1'h0 ),
       .io_cp_resp_valid( FPU_io_cp_resp_valid ),
       .io_cp_resp_bits_data( FPU_io_cp_resp_bits_data )
       //.io_cp_resp_bits_exc(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign FPU.io_cp_req_bits_cmd = {1{$random}};
    assign FPU.io_cp_req_bits_ldst = {1{$random}};
    assign FPU.io_cp_req_bits_wen = {1{$random}};
    assign FPU.io_cp_req_bits_ren1 = {1{$random}};
    assign FPU.io_cp_req_bits_ren2 = {1{$random}};
    assign FPU.io_cp_req_bits_ren3 = {1{$random}};
    assign FPU.io_cp_req_bits_swap12 = {1{$random}};
    assign FPU.io_cp_req_bits_swap23 = {1{$random}};
    assign FPU.io_cp_req_bits_single = {1{$random}};
    assign FPU.io_cp_req_bits_fromint = {1{$random}};
    assign FPU.io_cp_req_bits_toint = {1{$random}};
    assign FPU.io_cp_req_bits_fastpipe = {1{$random}};
    assign FPU.io_cp_req_bits_fma = {1{$random}};
    assign FPU.io_cp_req_bits_div = {1{$random}};
    assign FPU.io_cp_req_bits_sqrt = {1{$random}};
    assign FPU.io_cp_req_bits_round = {1{$random}};
    assign FPU.io_cp_req_bits_wflags = {1{$random}};
    assign FPU.io_cp_req_bits_rm = {1{$random}};
    assign FPU.io_cp_req_bits_typ = {1{$random}};
    assign FPU.io_cp_req_bits_in1 = {3{$random}};
    assign FPU.io_cp_req_bits_in2 = {3{$random}};
    assign FPU.io_cp_req_bits_in3 = {3{$random}};
// synthesis translate_on
`endif
  ClientTileLinkIOArbiter ClientTileLinkIOArbiter(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( ClientTileLinkIOArbiter_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( SampleAccel_io_autl_acquire_valid ),
       //.io_in_1_acquire_bits_addr_block(  )
       //.io_in_1_acquire_bits_client_xact_id(  )
       //.io_in_1_acquire_bits_addr_beat(  )
       //.io_in_1_acquire_bits_is_builtin_type(  )
       //.io_in_1_acquire_bits_a_type(  )
       //.io_in_1_acquire_bits_union(  )
       //.io_in_1_acquire_bits_data(  )
       .io_in_1_grant_ready( SampleAccel_io_autl_grant_ready ),
       .io_in_1_grant_valid( ClientTileLinkIOArbiter_io_in_1_grant_valid ),
       .io_in_1_grant_bits_addr_beat( ClientTileLinkIOArbiter_io_in_1_grant_bits_addr_beat ),
       .io_in_1_grant_bits_client_xact_id( ClientTileLinkIOArbiter_io_in_1_grant_bits_client_xact_id ),
       .io_in_1_grant_bits_manager_xact_id( ClientTileLinkIOArbiter_io_in_1_grant_bits_manager_xact_id ),
       .io_in_1_grant_bits_is_builtin_type( ClientTileLinkIOArbiter_io_in_1_grant_bits_is_builtin_type ),
       .io_in_1_grant_bits_g_type( ClientTileLinkIOArbiter_io_in_1_grant_bits_g_type ),
       .io_in_1_grant_bits_data( ClientTileLinkIOArbiter_io_in_1_grant_bits_data ),
       //.io_in_1_probe_ready(  )
       //.io_in_1_probe_valid(  )
       //.io_in_1_probe_bits_addr_block(  )
       //.io_in_1_probe_bits_p_type(  )
       //.io_in_1_release_ready(  )
       //.io_in_1_release_valid(  )
       //.io_in_1_release_bits_addr_beat(  )
       //.io_in_1_release_bits_addr_block(  )
       //.io_in_1_release_bits_client_xact_id(  )
       //.io_in_1_release_bits_voluntary(  )
       //.io_in_1_release_bits_r_type(  )
       //.io_in_1_release_bits_data(  )
       .io_in_0_acquire_ready( ClientTileLinkIOArbiter_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( icache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_in_0_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_in_0_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_in_0_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_in_0_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_in_0_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_in_0_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_in_0_grant_ready( icache_io_mem_grant_ready ),
       .io_in_0_grant_valid( ClientTileLinkIOArbiter_io_in_0_grant_valid ),
       .io_in_0_grant_bits_addr_beat( ClientTileLinkIOArbiter_io_in_0_grant_bits_addr_beat ),
       .io_in_0_grant_bits_client_xact_id( ClientTileLinkIOArbiter_io_in_0_grant_bits_client_xact_id ),
       .io_in_0_grant_bits_manager_xact_id( ClientTileLinkIOArbiter_io_in_0_grant_bits_manager_xact_id ),
       .io_in_0_grant_bits_is_builtin_type( ClientTileLinkIOArbiter_io_in_0_grant_bits_is_builtin_type ),
       .io_in_0_grant_bits_g_type( ClientTileLinkIOArbiter_io_in_0_grant_bits_g_type ),
       .io_in_0_grant_bits_data( ClientTileLinkIOArbiter_io_in_0_grant_bits_data ),
       //.io_in_0_probe_ready(  )
       //.io_in_0_probe_valid(  )
       //.io_in_0_probe_bits_addr_block(  )
       //.io_in_0_probe_bits_p_type(  )
       //.io_in_0_release_ready(  )
       //.io_in_0_release_valid(  )
       //.io_in_0_release_bits_addr_beat(  )
       //.io_in_0_release_bits_addr_block(  )
       //.io_in_0_release_bits_client_xact_id(  )
       //.io_in_0_release_bits_voluntary(  )
       //.io_in_0_release_bits_r_type(  )
       //.io_in_0_release_bits_data(  )
       .io_out_acquire_ready( io_uncached_0_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOArbiter_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOArbiter_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOArbiter_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOArbiter_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOArbiter_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOArbiter_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOArbiter_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOArbiter_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOArbiter_io_out_grant_ready ),
       .io_out_grant_valid( io_uncached_0_grant_valid ),
       .io_out_grant_bits_addr_beat( io_uncached_0_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( io_uncached_0_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( io_uncached_0_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( io_uncached_0_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( io_uncached_0_grant_bits_g_type ),
       .io_out_grant_bits_data( io_uncached_0_grant_bits_data )
       //.io_out_probe_ready(  )
       //.io_out_probe_valid(  )
       //.io_out_probe_bits_addr_block(  )
       //.io_out_probe_bits_p_type(  )
       //.io_out_release_ready(  )
       //.io_out_release_valid(  )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_addr_block = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_addr_beat = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_is_builtin_type = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_a_type = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_union = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_acquire_bits_data = {4{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_probe_ready = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_valid = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_addr_beat = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_addr_block = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_voluntary = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_r_type = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_1_release_bits_data = {4{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_probe_ready = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_valid = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_addr_beat = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_addr_block = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_voluntary = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_r_type = {1{$random}};
    assign ClientTileLinkIOArbiter.io_in_0_release_bits_data = {4{$random}};
    assign ClientTileLinkIOArbiter.io_out_probe_valid = {1{$random}};
    assign ClientTileLinkIOArbiter.io_out_probe_bits_addr_block = {1{$random}};
    assign ClientTileLinkIOArbiter.io_out_probe_bits_p_type = {1{$random}};
    assign ClientTileLinkIOArbiter.io_out_release_ready = {1{$random}};
// synthesis translate_on
`endif
  RRArbiter_0 RRArbiter(.clk(clk), .reset(reset),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( Queue_io_deq_valid ),
       .io_in_0_bits_rd( Queue_io_deq_bits_rd ),
       .io_in_0_bits_data( Queue_io_deq_bits_data ),
       .io_out_ready( core_io_rocc_resp_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_rd( RRArbiter_io_out_bits_rd ),
       .io_out_bits_data( RRArbiter_io_out_bits_data )
       //.io_chosen(  )
  );
  RoccCommandRouter RoccCommandRouter(.clk(clk), .reset(reset),
       .io_in_ready( RoccCommandRouter_io_in_ready ),
       .io_in_valid( core_io_rocc_cmd_valid ),
       .io_in_bits_inst_funct( core_io_rocc_cmd_bits_inst_funct ),
       .io_in_bits_inst_rs2( core_io_rocc_cmd_bits_inst_rs2 ),
       .io_in_bits_inst_rs1( core_io_rocc_cmd_bits_inst_rs1 ),
       .io_in_bits_inst_xd( core_io_rocc_cmd_bits_inst_xd ),
       .io_in_bits_inst_xs1( core_io_rocc_cmd_bits_inst_xs1 ),
       .io_in_bits_inst_xs2( core_io_rocc_cmd_bits_inst_xs2 ),
       .io_in_bits_inst_rd( core_io_rocc_cmd_bits_inst_rd ),
       .io_in_bits_inst_opcode( core_io_rocc_cmd_bits_inst_opcode ),
       .io_in_bits_rs1( core_io_rocc_cmd_bits_rs1 ),
       .io_in_bits_rs2( core_io_rocc_cmd_bits_rs2 ),
       .io_out_0_ready( SampleAccel_io_cmd_ready ),
       .io_out_0_valid( RoccCommandRouter_io_out_0_valid ),
       .io_out_0_bits_inst_funct( RoccCommandRouter_io_out_0_bits_inst_funct ),
       .io_out_0_bits_inst_rs2( RoccCommandRouter_io_out_0_bits_inst_rs2 ),
       .io_out_0_bits_inst_rs1( RoccCommandRouter_io_out_0_bits_inst_rs1 ),
       .io_out_0_bits_inst_xd( RoccCommandRouter_io_out_0_bits_inst_xd ),
       .io_out_0_bits_inst_xs1( RoccCommandRouter_io_out_0_bits_inst_xs1 ),
       .io_out_0_bits_inst_xs2( RoccCommandRouter_io_out_0_bits_inst_xs2 ),
       .io_out_0_bits_inst_rd( RoccCommandRouter_io_out_0_bits_inst_rd ),
       .io_out_0_bits_inst_opcode( RoccCommandRouter_io_out_0_bits_inst_opcode ),
       .io_out_0_bits_rs1( RoccCommandRouter_io_out_0_bits_rs1 ),
       .io_out_0_bits_rs2( RoccCommandRouter_io_out_0_bits_rs2 ),
       .io_busy( RoccCommandRouter_io_busy )
  );
  
  always @ (posedge clk) begin
    //$display(RoccCommandRouter_io_out_0_valid);
    if (RoccCommandRouter_io_out_0_valid) begin
      $display("1");
    end
  end
  
  mem_Accel_B SampleAccel(.clk(clk), .rst(reset),
       .cmd_rdy( SampleAccel_io_cmd_ready ),
       .cmd_vld( RoccCommandRouter_io_out_0_valid ),
       .cmd({
                  RoccCommandRouter_io_out_0_bits_rs2,
                  RoccCommandRouter_io_out_0_bits_rs1,
                  RoccCommandRouter_io_out_0_bits_inst_opcode,
                  RoccCommandRouter_io_out_0_bits_inst_rd,
                  RoccCommandRouter_io_out_0_bits_inst_xs2,
                  RoccCommandRouter_io_out_0_bits_inst_xs1,
                  RoccCommandRouter_io_out_0_bits_inst_xd,
                  RoccCommandRouter_io_out_0_bits_inst_rs1,
                  RoccCommandRouter_io_out_0_bits_inst_rs2,
                  RoccCommandRouter_io_out_0_bits_inst_funct
                  }),
       .resp_rdy( Queue_io_enq_ready ),
       .resp_vld( SampleAccel_io_resp_valid ),
       .resp({
                   SampleAccel_io_resp_bits_data,
                   SampleAccel_io_resp_bits_rd,
                   SampleAccel_io_mem_req_valid,
                   SampleAccel_io_autl_acquire_valid,
                   ClientTileLinkIOArbiter_io_in_1_acquire_ready,
                   SampleAccel_io_interrupt,
                   SampleAccel_io_busy
                   }),
       .mem_req_rdy( SimpleHellaCacheIF_io_requestor_req_ready ),
       .mem_req_vld( SimpleHellaCacheIF_io_requestor_req_valid ),
       .mem_req({
                      SimpleHellaCacheIF_io_requestor_req_addr,
                      SimpleHellaCacheIF_io_requestor_req_tag,
                      SimpleHellaCacheIF_io_requestor_req_cmd,
                      SimpleHellaCacheIF_io_requestor_req_typ, 
                      SimpleHellaCacheIF_io_requestor_req_kill, 
                      SimpleHellaCacheIF_io_requestor_req_phys, 
                      SimpleHellaCacheIF_io_requestor_req_data
                     }),
       //.io_mem_resp_V_ap_ack( ),
       .mem_resp_vld( SimpleHellaCacheIF_io_requestor_resp_valid ),
       .mem_resp({
                        SimpleHellaCacheIF_io_requestor_resp_bits_addr,
                        SimpleHellaCacheIF_io_requestor_resp_bits_tag,
                        SimpleHellaCacheIF_io_requestor_resp_bits_cmd,
                        SimpleHellaCacheIF_io_requestor_resp_bits_typ,
                        SimpleHellaCacheIF_io_requestor_resp_bits_data,
                        SimpleHellaCacheIF_io_requestor_resp_bits_nack,
                        SimpleHellaCacheIF_io_requestor_resp_bits_replay,
                        SimpleHellaCacheIF_io_requestor_resp_bits_has_data,
                        SimpleHellaCacheIF_io_requestor_resp_bits_data_word_bypass,
                        SimpleHellaCacheIF_io_requestor_resp_bits_store_data 
                     })
  );
  
  /*
  reg toggle;
  
  always @ (posedge clk) begin
    if (reset) begin
      toggle <= 1'b0;
    end
    if (RoccCommandRouter_io_out_0_valid) begin
      toggle <= 1'b1;
      $display("~~~~~");
      $display("RoccCommandRouter_io_out_0_valid:");
      $display(RoccCommandRouter_io_out_0_valid);
      $display("------");
      $display("rst:");
      $display(SampleAccel.rst);
      $display("state_reg:");
      $display(SampleAccel.state_reg);
      $display("next_state:");
      $display(SampleAccel.next_state);
      $display("cmd_vld:");
      $display(SampleAccel.cmd_vld);
      $display("cmd_rdy:");
      $display(SampleAccel.cmd_rdy);
      $display("cmd_go:");
      $display(SampleAccel.cmd_go);
      $display("resp_vld:");
      $display(SampleAccel.resp_vld);
      $display("resp_rdy:");
      $display(SampleAccel.resp_rdy);
      $display("resp_go:");
      $display(SampleAccel.resp_go);
      $display("------");
      $display("rs1_data:");
      $display(SampleAccel.cmd_rs1_data);
      $display("rs2_data:");
      $display(SampleAccel.cmd_rs2_data);
      $display("adder_out:");
      $display(SampleAccel.adder_out);
      $display("resp_data:");
      $display(SampleAccel.resp_data);
      $display("------");
      $display("cmd_inst_rd:");
      $display(SampleAccel.cmd_inst_rd);
      $display("resp_rd:");
      $display(SampleAccel.resp_rd);
      $display("------");
    end
    if (toggle) begin
      toggle <= 1'b0;
      $display("~~~~~");
      $display("RoccCommandRouter_io_out_0_valid:");
      $display(RoccCommandRouter_io_out_0_valid);
      $display("------");
      $display("rst:");
      $display(SampleAccel.rst);
      $display("state_reg:");
      $display(SampleAccel.state_reg);
      $display("next_state:");
      $display(SampleAccel.next_state);
      $display("cmd_vld:");
      $display(SampleAccel.cmd_vld);
      $display("cmd_rdy:");
      $display(SampleAccel.cmd_rdy);
      $display("cmd_go:");
      $display(SampleAccel.cmd_go);
      $display("resp_vld:");
      $display(SampleAccel.resp_vld);
      $display("resp_rdy:");
      $display(SampleAccel.resp_rdy);
      $display("resp_go:");
      $display(SampleAccel.resp_go);
      $display("------");
      $display("rs1_data:");
      $display(SampleAccel.cmd_rs1_data);
      $display("rs2_data:");
      $display(SampleAccel.cmd_rs2_data);
      $display("adder_out:");
      $display(SampleAccel.adder_out);
      $display("resp_data:");
      $display(SampleAccel.resp_data);
      $display("------");
      $display("cmd_inst_rd:");
      $display(SampleAccel.cmd_inst_rd);
      $display("resp_rd:");
      $display(SampleAccel.resp_rd);
      $display("------");
    end
  end
  
  // Yangyi
  adder_Accel SampleAccel
  (
    .clk      ( clk ),
    .rst      ( reset ),
    .cmd      ({
                RoccCommandRouter_io_out_0_bits_rs2,
                RoccCommandRouter_io_out_0_bits_rs1,
                RoccCommandRouter_io_out_0_bits_inst_opcode,
                RoccCommandRouter_io_out_0_bits_inst_rd,
                RoccCommandRouter_io_out_0_bits_inst_xs2,
                RoccCommandRouter_io_out_0_bits_inst_xs1,
                RoccCommandRouter_io_out_0_bits_inst_xd,
                RoccCommandRouter_io_out_0_bits_inst_rs1,
                RoccCommandRouter_io_out_0_bits_inst_rs2,
                RoccCommandRouter_io_out_0_bits_inst_funct
              }),
    .cmd_vld  ( RoccCommandRouter_io_out_0_valid ),
    .cmd_rdy  ( SampleAccel_io_cmd_ready ),
    .resp     ({
                SampleAccel_io_resp_bits_data,
                SampleAccel_io_resp_bits_rd,
                SampleAccel_io_mem_req_valid,
                SampleAccel_io_autl_acquire_valid,
                ClientTileLinkIOArbiter_io_in_1_acquire_ready,
                SampleAccel_io_interrupt,
                SampleAccel_io_busy
              }),
    .resp_vld ( SampleAccel_io_resp_valid ),
    .resp_rdy ( Queue_io_enq_ready )
  );
  */
  /*
  //gai
  gcd SampleAccel(.ap_clk(clk), .ap_rst(reset),
       .io_cmd_V_ap_ack( SampleAccel_io_cmd_ready ),
       .io_cmd_V_ap_vld( RoccCommandRouter_io_out_0_valid ),
       .io_cmd_V({
                  RoccCommandRouter_io_out_0_bits_rs2,
                  RoccCommandRouter_io_out_0_bits_rs1,
                  RoccCommandRouter_io_out_0_bits_inst_opcode,
                  RoccCommandRouter_io_out_0_bits_inst_rd,
                  RoccCommandRouter_io_out_0_bits_inst_xs2,
                  RoccCommandRouter_io_out_0_bits_inst_xs1,
                  RoccCommandRouter_io_out_0_bits_inst_xd,
                  RoccCommandRouter_io_out_0_bits_inst_rs1,
                  RoccCommandRouter_io_out_0_bits_inst_rs2,
                  RoccCommandRouter_io_out_0_bits_inst_funct
                  }),
       //.io_cmd_V[6:0]( RoccCommandRouter_io_out_0_bits_inst_funct ),
       //.io_cmd_V[11:7]( RoccCommandRouter_io_out_0_bits_inst_rs2 ),
       //.io_cmd_V[16:12]( RoccCommandRouter_io_out_0_bits_inst_rs1 ),
       //.io_cmd_V[17]( RoccCommandRouter_io_out_0_bits_inst_xd ),
       //.io_cmd_V[18]( RoccCommandRouter_io_out_0_bits_inst_xs1 ),
       //.io_cmd_V[19]( RoccCommandRouter_io_out_0_bits_inst_xs2 ),
       //.io_cmd_V[24:20]( RoccCommandRouter_io_out_0_bits_inst_rd ),
       //.io_cmd_V[31:25]( RoccCommandRouter_io_out_0_bits_inst_opcode ),
       //.io_cmd_V[95:32]( RoccCommandRouter_io_out_0_bits_rs1 ),
       //.io_cmd_V[159:96]( RoccCommandRouter_io_out_0_bits_rs2 ),
       .io_resp_V_ap_ack( Queue_io_enq_ready ),
       .io_resp_V_ap_vld( SampleAccel_io_resp_valid ),
       .io_resp_V({
                   SampleAccel_io_resp_bits_data,
                   SampleAccel_io_resp_bits_rd,
                   SampleAccel_io_mem_req_valid,
                   SampleAccel_io_autl_acquire_valid,
                   ClientTileLinkIOArbiter_io_in_1_acquire_ready,
                   SampleAccel_io_interrupt,
                   SampleAccel_io_busy
                   })
       //.io_resp_V[0]( SampleAccel_io_busy ),
       //.io_resp_V[1]( SampleAccel_io_interrupt ),
       //.io_resp_V[2]( ClientTileLinkIOArbiter_io_in_1_acquire_ready ),
       //.io_resp_V[3]( SampleAccel_io_autl_acquire_valid ),
       //.io_resp_V[4]( SampleAccel_io_mem_req_valid ),
       //.io_resp_V[9:5]( SampleAccel_io_resp_bits_rd ),
       //.io_resp_V[73:10]( SampleAccel_io_resp_bits_data )
       //.io_mem_req_ready( SimpleHellaCacheIF_io_requestor_req_ready ),
       //.io_mem_req_bits_addr(  )
       //.io_mem_req_bits_tag(  )
       //.io_mem_req_bits_cmd(  )
       //.io_mem_req_bits_typ(  )
       //.io_mem_req_bits_kill(  )
       //.io_mem_req_bits_phys( SampleAccel_io_mem_req_bits_phys ),
       //.io_mem_req_bits_data(  )
       //.io_mem_resp_valid( SimpleHellaCacheIF_io_requestor_resp_valid ),
       //.io_mem_resp_bits_addr( SimpleHellaCacheIF_io_requestor_resp_bits_addr ),
       //.io_mem_resp_bits_tag( SimpleHellaCacheIF_io_requestor_resp_bits_tag ),
       //.io_mem_resp_bits_cmd( SimpleHellaCacheIF_io_requestor_resp_bits_cmd ),
       //.io_mem_resp_bits_typ( SimpleHellaCacheIF_io_requestor_resp_bits_typ ),
       //.io_mem_resp_bits_data( SimpleHellaCacheIF_io_requestor_resp_bits_data ),
       //.io_mem_resp_bits_nack( SimpleHellaCacheIF_io_requestor_resp_bits_nack ),
       //.io_mem_resp_bits_replay( SimpleHellaCacheIF_io_requestor_resp_bits_replay ),
       //.io_mem_resp_bits_has_data( SimpleHellaCacheIF_io_requestor_resp_bits_has_data ),
       //.io_mem_resp_bits_data_word_bypass( SimpleHellaCacheIF_io_requestor_resp_bits_data_word_bypass ),
       //.io_mem_resp_bits_store_data( SimpleHellaCacheIF_io_requestor_resp_bits_store_data ),
       //.io_mem_replay_next_valid(  )
       //.io_mem_replay_next_bits(  )
       //.io_mem_xcpt_ma_ld(  )
       //.io_mem_xcpt_ma_st(  )
       //.io_mem_xcpt_pf_ld(  )
       //.io_mem_xcpt_pf_st(  )
       //.io_mem_invalidate_lr(  )
       //.io_mem_ordered(  )
       //.io_s( core_io_rocc_s ),
       //.io_autl_acquire_bits_addr_block(  )
       //.io_autl_acquire_bits_client_xact_id(  )
       //.io_autl_acquire_bits_addr_beat(  )
       //.io_autl_acquire_bits_is_builtin_type(  )
       //.io_autl_acquire_bits_a_type(  )
       //.io_autl_acquire_bits_union(  )
       //.io_autl_acquire_bits_data(  )
       //.io_autl_grant_ready( SampleAccel_io_autl_grant_ready ),
       //.io_autl_grant_valid( ClientTileLinkIOArbiter_io_in_1_grant_valid ),
       //.io_autl_grant_bits_addr_beat( ClientTileLinkIOArbiter_io_in_1_grant_bits_addr_beat ),
       //.io_autl_grant_bits_client_xact_id( ClientTileLinkIOArbiter_io_in_1_grant_bits_client_xact_id ),
       //.io_autl_grant_bits_manager_xact_id( ClientTileLinkIOArbiter_io_in_1_grant_bits_manager_xact_id ),
       //.io_autl_grant_bits_is_builtin_type( ClientTileLinkIOArbiter_io_in_1_grant_bits_is_builtin_type ),
       //.io_autl_grant_bits_g_type( ClientTileLinkIOArbiter_io_in_1_grant_bits_g_type ),
       //.io_autl_grant_bits_data( ClientTileLinkIOArbiter_io_in_1_grant_bits_data ),
       //.io_fpu_req_ready(  )
       //.io_fpu_req_valid(  )
       //.io_fpu_req_bits_cmd(  )
       //.io_fpu_req_bits_ldst(  )
       //.io_fpu_req_bits_wen(  )
       //.io_fpu_req_bits_ren1(  )
       //.io_fpu_req_bits_ren2(  )
       //.io_fpu_req_bits_ren3(  )
       //.io_fpu_req_bits_swap12(  )
       //.io_fpu_req_bits_swap23(  )
       //.io_fpu_req_bits_single(  )
       //.io_fpu_req_bits_fromint(  )
       //.io_fpu_req_bits_toint(  )
       //.io_fpu_req_bits_fastpipe(  )
       //.io_fpu_req_bits_fma(  )
       //.io_fpu_req_bits_div(  )
       //.io_fpu_req_bits_sqrt(  )
       //.io_fpu_req_bits_round(  )
       //.io_fpu_req_bits_wflags(  )
       //.io_fpu_req_bits_rm(  )
       //.io_fpu_req_bits_typ(  )
       //.io_fpu_req_bits_in1(  )
       //.io_fpu_req_bits_in2(  )
       //.io_fpu_req_bits_in3(  )
       //.io_fpu_resp_ready(  )
       //.io_fpu_resp_valid(  )
       //.io_fpu_resp_bits_data(  )
       //.io_fpu_resp_bits_exc(  )
       //.io_exception( core_io_rocc_exception ),
       //.io_csr_waddr(  )
       //.io_csr_wdata(  )
       //.io_csr_wen(  )
       //.io_host_id( io_host_id )
  );
  */
  SimpleHellaCacheIF SimpleHellaCacheIF(.clk(clk), .reset(reset),
       .io_requestor_req_ready( SimpleHellaCacheIF_io_requestor_req_ready ),
       .io_requestor_req_valid( SampleAccel_io_mem_req_valid ),
       .io_requestor_req_bits_addr( SimpleHellaCacheIF_io_requestor_req_addr ),
       .io_requestor_req_bits_tag( SimpleHellaCacheIF_io_requestor_req_tag ),
       .io_requestor_req_bits_cmd( SimpleHellaCacheIF_io_requestor_req_cmd ),
       .io_requestor_req_bits_typ( SimpleHellaCacheIF_io_requestor_req_typ ),
       .io_requestor_req_bits_kill( SimpleHellaCacheIF_io_requestor_req_kill ),
       .io_requestor_req_bits_phys( SampleAccel_io_mem_req_bits_phys ),
       .io_requestor_req_bits_data( SimpleHellaCacheIF_io_requestor_req_data ),
       .io_requestor_resp_valid( SimpleHellaCacheIF_io_requestor_resp_valid ),
       .io_requestor_resp_bits_addr( SimpleHellaCacheIF_io_requestor_resp_bits_addr ),
       .io_requestor_resp_bits_tag( SimpleHellaCacheIF_io_requestor_resp_bits_tag ),
       .io_requestor_resp_bits_cmd( SimpleHellaCacheIF_io_requestor_resp_bits_cmd ),
       .io_requestor_resp_bits_typ( SimpleHellaCacheIF_io_requestor_resp_bits_typ ),
       .io_requestor_resp_bits_data( SimpleHellaCacheIF_io_requestor_resp_bits_data ),
       .io_requestor_resp_bits_nack( SimpleHellaCacheIF_io_requestor_resp_bits_nack ),
       .io_requestor_resp_bits_replay( SimpleHellaCacheIF_io_requestor_resp_bits_replay ),
       .io_requestor_resp_bits_has_data( SimpleHellaCacheIF_io_requestor_resp_bits_has_data ),
       .io_requestor_resp_bits_data_word_bypass( SimpleHellaCacheIF_io_requestor_resp_bits_data_word_bypass ),
       .io_requestor_resp_bits_store_data( SimpleHellaCacheIF_io_requestor_resp_bits_store_data ),
       //.io_requestor_replay_next_valid(  )
       //.io_requestor_replay_next_bits(  )
       //.io_requestor_xcpt_ma_ld(  )
       //.io_requestor_xcpt_ma_st(  )
       //.io_requestor_xcpt_pf_ld(  )
       //.io_requestor_xcpt_pf_st(  )
       //.io_requestor_invalidate_lr(  )
       //.io_requestor_ordered(  )
       .io_cache_req_ready( dcArb_io_requestor_2_req_ready ),
       .io_cache_req_valid( SimpleHellaCacheIF_io_cache_req_valid ),
       .io_cache_req_bits_addr( SimpleHellaCacheIF_io_cache_req_bits_addr ),
       .io_cache_req_bits_tag( SimpleHellaCacheIF_io_cache_req_bits_tag ),
       .io_cache_req_bits_cmd( SimpleHellaCacheIF_io_cache_req_bits_cmd ),
       .io_cache_req_bits_typ( SimpleHellaCacheIF_io_cache_req_bits_typ ),
       .io_cache_req_bits_kill( SimpleHellaCacheIF_io_cache_req_bits_kill ),
       .io_cache_req_bits_phys( SimpleHellaCacheIF_io_cache_req_bits_phys ),
       .io_cache_req_bits_data( SimpleHellaCacheIF_io_cache_req_bits_data ),
       .io_cache_resp_valid( dcArb_io_requestor_2_resp_valid ),
       .io_cache_resp_bits_addr( dcArb_io_requestor_2_resp_bits_addr ),
       .io_cache_resp_bits_tag( dcArb_io_requestor_2_resp_bits_tag ),
       .io_cache_resp_bits_cmd( dcArb_io_requestor_2_resp_bits_cmd ),
       .io_cache_resp_bits_typ( dcArb_io_requestor_2_resp_bits_typ ),
       .io_cache_resp_bits_data( dcArb_io_requestor_2_resp_bits_data ),
       .io_cache_resp_bits_nack( dcArb_io_requestor_2_resp_bits_nack ),
       .io_cache_resp_bits_replay( dcArb_io_requestor_2_resp_bits_replay ),
       .io_cache_resp_bits_has_data( dcArb_io_requestor_2_resp_bits_has_data ),
       .io_cache_resp_bits_data_word_bypass( dcArb_io_requestor_2_resp_bits_data_word_bypass ),
       .io_cache_resp_bits_store_data( dcArb_io_requestor_2_resp_bits_store_data ),
       .io_cache_replay_next_valid( dcArb_io_requestor_2_replay_next_valid ),
       .io_cache_replay_next_bits( dcArb_io_requestor_2_replay_next_bits ),
       .io_cache_xcpt_ma_ld( dcArb_io_requestor_2_xcpt_ma_ld ),
       .io_cache_xcpt_ma_st( dcArb_io_requestor_2_xcpt_ma_st ),
       .io_cache_xcpt_pf_ld( dcArb_io_requestor_2_xcpt_pf_ld ),
       .io_cache_xcpt_pf_st( dcArb_io_requestor_2_xcpt_pf_st ),
       //.io_cache_invalidate_lr(  )
       .io_cache_ordered( dcArb_io_requestor_2_ordered )
  );
//`ifndef SYNTHESIS
//// synthesis translate_off
//    assign SimpleHellaCacheIF.io_requestor_req_bits_addr = {2{$random}};
//    assign SimpleHellaCacheIF.io_requestor_req_bits_tag = {1{$random}};
//    assign SimpleHellaCacheIF.io_requestor_req_bits_cmd = {1{$random}};
//    assign SimpleHellaCacheIF.io_requestor_req_bits_typ = {1{$random}};
//    assign SimpleHellaCacheIF.io_requestor_req_bits_kill = {1{$random}};
//    assign SimpleHellaCacheIF.io_requestor_req_bits_data = {2{$random}};
//// synthesis translate_on
//`endif
  Queue_6 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( SampleAccel_io_resp_valid ),
       .io_enq_bits_rd( SampleAccel_io_resp_bits_rd ),
       .io_enq_bits_data( SampleAccel_io_resp_bits_data ),
       .io_deq_ready( RRArbiter_io_in_0_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_rd( Queue_io_deq_bits_rd ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [11:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[11:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[76:0] T11;
  reg [76:0] ram [1:0];
  wire[76:0] T12;
  wire[76:0] T13;
  wire[76:0] T14;
  wire[75:0] T15;
  wire[11:0] T16;
  wire T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rw, T15};
  assign T15 = {io_enq_bits_addr, io_enq_bits_data};
  assign io_deq_bits_addr = T16;
  assign T16 = T11[7'h4b:7'h40];
  assign io_deq_bits_rw = T17;
  assign T17 = T11[7'h4c];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[63:0] T10;
  reg [63:0] ram [1:0];
  wire[63:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    output io_mem_backup_ctrl_out_valid,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[5:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [5:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[5:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [5:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    input  init
);

  reg  R0;
  reg  R1;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire Queue_io_deq_bits_rw;
  wire[11:0] Queue_io_deq_bits_addr;
  wire[63:0] Queue_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[31:0] Queue_2_io_deq_bits_addr;
  wire[7:0] Queue_2_io_deq_bits_len;
  wire[2:0] Queue_2_io_deq_bits_size;
  wire[1:0] Queue_2_io_deq_bits_burst;
  wire Queue_2_io_deq_bits_lock;
  wire[2:0] Queue_2_io_deq_bits_prot;
  wire[3:0] Queue_2_io_deq_bits_qos;
  wire[3:0] Queue_2_io_deq_bits_region;
  wire[5:0] Queue_2_io_deq_bits_id;
  wire Queue_2_io_deq_bits_user;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[31:0] Queue_3_io_deq_bits_addr;
  wire[7:0] Queue_3_io_deq_bits_len;
  wire[2:0] Queue_3_io_deq_bits_size;
  wire[1:0] Queue_3_io_deq_bits_burst;
  wire Queue_3_io_deq_bits_lock;
  wire[2:0] Queue_3_io_deq_bits_prot;
  wire[3:0] Queue_3_io_deq_bits_qos;
  wire[3:0] Queue_3_io_deq_bits_region;
  wire[5:0] Queue_3_io_deq_bits_id;
  wire Queue_3_io_deq_bits_user;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[63:0] Queue_4_io_deq_bits_data;
  wire Queue_4_io_deq_bits_last;
  wire[7:0] Queue_4_io_deq_bits_strb;
  wire Queue_4_io_deq_bits_user;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_resp;
  wire[63:0] Queue_5_io_deq_bits_data;
  wire Queue_5_io_deq_bits_last;
  wire[5:0] Queue_5_io_deq_bits_id;
  wire Queue_5_io_deq_bits_user;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_resp;
  wire[5:0] Queue_6_io_deq_bits_id;
  wire Queue_6_io_deq_bits_user;
  wire RocketTile_io_cached_0_acquire_valid;
  wire[25:0] RocketTile_io_cached_0_acquire_bits_addr_block;
  wire[5:0] RocketTile_io_cached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_cached_0_acquire_bits_addr_beat;
  wire RocketTile_io_cached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_cached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_cached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_cached_0_acquire_bits_data;
  wire RocketTile_io_cached_0_grant_ready;
  wire RocketTile_io_cached_0_probe_ready;
  wire RocketTile_io_cached_0_release_valid;
  wire[1:0] RocketTile_io_cached_0_release_bits_addr_beat;
  wire[25:0] RocketTile_io_cached_0_release_bits_addr_block;
  wire[5:0] RocketTile_io_cached_0_release_bits_client_xact_id;
  wire RocketTile_io_cached_0_release_bits_voluntary;
  wire[2:0] RocketTile_io_cached_0_release_bits_r_type;
  wire[127:0] RocketTile_io_cached_0_release_bits_data;
  wire RocketTile_io_uncached_0_acquire_valid;
  wire[25:0] RocketTile_io_uncached_0_acquire_bits_addr_block;
  wire[5:0] RocketTile_io_uncached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_uncached_0_acquire_bits_addr_beat;
  wire RocketTile_io_uncached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_uncached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_uncached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_uncached_0_acquire_bits_data;
  wire RocketTile_io_uncached_0_grant_ready;
  wire RocketTile_io_host_csr_req_ready;
  wire RocketTile_io_host_csr_resp_valid;
  wire[63:0] RocketTile_io_host_csr_resp_bits;
  wire RocketTile_io_host_debug_stats_csr;
  wire uncore_io_host_clk;
  wire uncore_io_host_clk_edge;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_csr;
  wire uncore_io_mem_0_aw_valid;
  wire[31:0] uncore_io_mem_0_aw_bits_addr;
  wire[7:0] uncore_io_mem_0_aw_bits_len;
  wire[2:0] uncore_io_mem_0_aw_bits_size;
  wire[1:0] uncore_io_mem_0_aw_bits_burst;
  wire uncore_io_mem_0_aw_bits_lock;
  wire[3:0] uncore_io_mem_0_aw_bits_cache;
  wire[2:0] uncore_io_mem_0_aw_bits_prot;
  wire[3:0] uncore_io_mem_0_aw_bits_qos;
  wire[3:0] uncore_io_mem_0_aw_bits_region;
  wire[5:0] uncore_io_mem_0_aw_bits_id;
  wire uncore_io_mem_0_aw_bits_user;
  wire uncore_io_mem_0_w_valid;
  wire[63:0] uncore_io_mem_0_w_bits_data;
  wire uncore_io_mem_0_w_bits_last;
  wire[7:0] uncore_io_mem_0_w_bits_strb;
  wire uncore_io_mem_0_w_bits_user;
  wire uncore_io_mem_0_b_ready;
  wire uncore_io_mem_0_ar_valid;
  wire[31:0] uncore_io_mem_0_ar_bits_addr;
  wire[7:0] uncore_io_mem_0_ar_bits_len;
  wire[2:0] uncore_io_mem_0_ar_bits_size;
  wire[1:0] uncore_io_mem_0_ar_bits_burst;
  wire uncore_io_mem_0_ar_bits_lock;
  wire[3:0] uncore_io_mem_0_ar_bits_cache;
  wire[2:0] uncore_io_mem_0_ar_bits_prot;
  wire[3:0] uncore_io_mem_0_ar_bits_qos;
  wire[3:0] uncore_io_mem_0_ar_bits_region;
  wire[5:0] uncore_io_mem_0_ar_bits_id;
  wire uncore_io_mem_0_ar_bits_user;
  wire uncore_io_mem_0_r_ready;
  wire uncore_io_tiles_cached_0_acquire_ready;
  wire uncore_io_tiles_cached_0_grant_valid;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire[5:0] uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire uncore_io_tiles_cached_0_probe_valid;
  wire[25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire uncore_io_tiles_cached_0_release_ready;
  wire uncore_io_tiles_uncached_0_acquire_ready;
  wire uncore_io_tiles_uncached_0_grant_valid;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[5:0] uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_csr_req_valid;
  wire uncore_io_htif_0_csr_req_bits_rw;
  wire[11:0] uncore_io_htif_0_csr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_csr_req_bits_data;
  wire uncore_io_htif_0_csr_resp_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_0_r_ready = Queue_5_io_enq_ready;
  assign io_mem_0_ar_bits_user = Queue_2_io_deq_bits_user;
  assign io_mem_0_ar_bits_id = Queue_2_io_deq_bits_id;
  assign io_mem_0_ar_bits_region = Queue_2_io_deq_bits_region;
  assign io_mem_0_ar_bits_qos = Queue_2_io_deq_bits_qos;
  assign io_mem_0_ar_bits_prot = Queue_2_io_deq_bits_prot;
  assign io_mem_0_ar_bits_cache = 4'h3;
  assign io_mem_0_ar_bits_lock = Queue_2_io_deq_bits_lock;
  assign io_mem_0_ar_bits_burst = Queue_2_io_deq_bits_burst;
  assign io_mem_0_ar_bits_size = Queue_2_io_deq_bits_size;
  assign io_mem_0_ar_bits_len = Queue_2_io_deq_bits_len;
  assign io_mem_0_ar_bits_addr = Queue_2_io_deq_bits_addr;
  assign io_mem_0_ar_valid = Queue_2_io_deq_valid;
  assign io_mem_0_b_ready = Queue_6_io_enq_ready;
  assign io_mem_0_w_bits_user = Queue_4_io_deq_bits_user;
  assign io_mem_0_w_bits_strb = Queue_4_io_deq_bits_strb;
  assign io_mem_0_w_bits_last = Queue_4_io_deq_bits_last;
  assign io_mem_0_w_bits_data = Queue_4_io_deq_bits_data;
  assign io_mem_0_w_valid = Queue_4_io_deq_valid;
  assign io_mem_0_aw_bits_user = Queue_3_io_deq_bits_user;
  assign io_mem_0_aw_bits_id = Queue_3_io_deq_bits_id;
  assign io_mem_0_aw_bits_region = Queue_3_io_deq_bits_region;
  assign io_mem_0_aw_bits_qos = Queue_3_io_deq_bits_qos;
  assign io_mem_0_aw_bits_prot = Queue_3_io_deq_bits_prot;
  assign io_mem_0_aw_bits_cache = 4'h3;
  assign io_mem_0_aw_bits_lock = Queue_3_io_deq_bits_lock;
  assign io_mem_0_aw_bits_burst = Queue_3_io_deq_bits_burst;
  assign io_mem_0_aw_bits_size = Queue_3_io_deq_bits_size;
  assign io_mem_0_aw_bits_len = Queue_3_io_deq_bits_len;
  assign io_mem_0_aw_bits_addr = Queue_3_io_deq_bits_addr;
  assign io_mem_0_aw_valid = Queue_3_io_deq_valid;
  assign io_host_debug_stats_csr = uncore_io_host_debug_stats_csr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  assign io_host_clk_edge = uncore_io_host_clk_edge;
  assign io_host_clk = uncore_io_host_clk;
  Uncore uncore(.clk(clk), .reset(reset),
       .io_host_clk( uncore_io_host_clk ),
       .io_host_clk_edge( uncore_io_host_clk_edge ),
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_csr( uncore_io_host_debug_stats_csr ),
       .io_mem_0_aw_ready( Queue_3_io_enq_ready ),
       .io_mem_0_aw_valid( uncore_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( Queue_4_io_enq_ready ),
       .io_mem_0_w_valid( uncore_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( uncore_io_mem_0_b_ready ),
       .io_mem_0_b_valid( Queue_6_io_deq_valid ),
       .io_mem_0_b_bits_resp( Queue_6_io_deq_bits_resp ),
       .io_mem_0_b_bits_id( Queue_6_io_deq_bits_id ),
       .io_mem_0_b_bits_user( Queue_6_io_deq_bits_user ),
       .io_mem_0_ar_ready( Queue_2_io_enq_ready ),
       .io_mem_0_ar_valid( uncore_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( uncore_io_mem_0_r_ready ),
       .io_mem_0_r_valid( Queue_5_io_deq_valid ),
       .io_mem_0_r_bits_resp( Queue_5_io_deq_bits_resp ),
       .io_mem_0_r_bits_data( Queue_5_io_deq_bits_data ),
       .io_mem_0_r_bits_last( Queue_5_io_deq_bits_last ),
       .io_mem_0_r_bits_id( Queue_5_io_deq_bits_id ),
       .io_mem_0_r_bits_user( Queue_5_io_deq_bits_user ),
       .io_tiles_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_csr_req_ready( Queue_io_enq_ready ),
       .io_htif_0_csr_req_valid( uncore_io_htif_0_csr_req_valid ),
       .io_htif_0_csr_req_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_htif_0_csr_req_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_htif_0_csr_req_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_htif_0_csr_resp_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_htif_0_csr_resp_valid( Queue_1_io_deq_valid ),
       .io_htif_0_csr_resp_bits( Queue_1_io_deq_bits ),
       .io_htif_0_debug_stats_csr( RocketTile_io_host_debug_stats_csr ),
       .io_mem_backup_ctrl_en( 1'h0 )
       //.io_mem_backup_ctrl_in_valid(  )
       //.io_mem_backup_ctrl_out_ready(  )
       //.io_mem_backup_ctrl_out_valid(  )
       //.io_mmio_aw_ready(  )
       //.io_mmio_aw_valid(  )
       //.io_mmio_aw_bits_addr(  )
       //.io_mmio_aw_bits_len(  )
       //.io_mmio_aw_bits_size(  )
       //.io_mmio_aw_bits_burst(  )
       //.io_mmio_aw_bits_lock(  )
       //.io_mmio_aw_bits_cache(  )
       //.io_mmio_aw_bits_prot(  )
       //.io_mmio_aw_bits_qos(  )
       //.io_mmio_aw_bits_region(  )
       //.io_mmio_aw_bits_id(  )
       //.io_mmio_aw_bits_user(  )
       //.io_mmio_w_ready(  )
       //.io_mmio_w_valid(  )
       //.io_mmio_w_bits_data(  )
       //.io_mmio_w_bits_last(  )
       //.io_mmio_w_bits_strb(  )
       //.io_mmio_w_bits_user(  )
       //.io_mmio_b_ready(  )
       //.io_mmio_b_valid(  )
       //.io_mmio_b_bits_resp(  )
       //.io_mmio_b_bits_id(  )
       //.io_mmio_b_bits_user(  )
       //.io_mmio_ar_ready(  )
       //.io_mmio_ar_valid(  )
       //.io_mmio_ar_bits_addr(  )
       //.io_mmio_ar_bits_len(  )
       //.io_mmio_ar_bits_size(  )
       //.io_mmio_ar_bits_burst(  )
       //.io_mmio_ar_bits_lock(  )
       //.io_mmio_ar_bits_cache(  )
       //.io_mmio_ar_bits_prot(  )
       //.io_mmio_ar_bits_qos(  )
       //.io_mmio_ar_bits_region(  )
       //.io_mmio_ar_bits_id(  )
       //.io_mmio_ar_bits_user(  )
       //.io_mmio_r_ready(  )
       //.io_mmio_r_valid(  )
       //.io_mmio_r_bits_resp(  )
       //.io_mmio_r_bits_data(  )
       //.io_mmio_r_bits_last(  )
       //.io_mmio_r_bits_id(  )
       //.io_mmio_r_bits_user(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign uncore.io_mem_backup_ctrl_in_valid = {1{$random}};
    assign uncore.io_mem_backup_ctrl_out_ready = {1{$random}};
// synthesis translate_on
`endif
  RocketTile RocketTile(.clk(clk), .reset(uncore_io_htif_0_reset),
       .io_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_csr_req_ready( RocketTile_io_host_csr_req_ready ),
       .io_host_csr_req_valid( Queue_io_deq_valid ),
       .io_host_csr_req_bits_rw( Queue_io_deq_bits_rw ),
       .io_host_csr_req_bits_addr( Queue_io_deq_bits_addr ),
       .io_host_csr_req_bits_data( Queue_io_deq_bits_data ),
       .io_host_csr_resp_ready( Queue_1_io_enq_ready ),
       .io_host_csr_resp_valid( RocketTile_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( RocketTile_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( RocketTile_io_host_debug_stats_csr ),
       //.io_dma_req_ready(  )
       //.io_dma_req_valid(  )
       //.io_dma_req_bits_xact_id(  )
       //.io_dma_req_bits_client_id(  )
       //.io_dma_req_bits_cmd(  )
       //.io_dma_req_bits_source(  )
       //.io_dma_req_bits_dest(  )
       //.io_dma_req_bits_length(  )
       //.io_dma_req_bits_size(  )
       //.io_dma_resp_ready(  )
       //.io_dma_resp_valid(  )
       //.io_dma_resp_bits_xact_id(  )
       //.io_dma_resp_bits_client_id(  )
       //.io_dma_resp_bits_status(  )
       .init( init )
  );
  Queue_0 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_csr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_csr_req_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_rw( Queue_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_csr_resp_valid ),
       .io_enq_bits( RocketTile_io_host_csr_resp_bits ),
       .io_deq_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_ar_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_deq_ready( io_mem_0_ar_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_addr( Queue_2_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_2_io_deq_bits_len ),
       .io_deq_bits_size( Queue_2_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_2_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_2_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_2_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_2_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_2_io_deq_bits_region ),
       .io_deq_bits_id( Queue_2_io_deq_bits_id ),
       .io_deq_bits_user( Queue_2_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_aw_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_deq_ready( io_mem_0_aw_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_addr( Queue_3_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_3_io_deq_bits_len ),
       .io_deq_bits_size( Queue_3_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_3_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_3_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_3_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_3_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_3_io_deq_bits_region ),
       .io_deq_bits_id( Queue_3_io_deq_bits_id ),
       .io_deq_bits_user( Queue_3_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_w_valid ),
       .io_enq_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_enq_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_enq_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_enq_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_deq_ready( io_mem_0_w_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_data( Queue_4_io_deq_bits_data ),
       .io_deq_bits_last( Queue_4_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_4_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( io_mem_0_r_valid ),
       .io_enq_bits_resp( io_mem_0_r_bits_resp ),
       .io_enq_bits_data( io_mem_0_r_bits_data ),
       .io_enq_bits_last( io_mem_0_r_bits_last ),
       .io_enq_bits_id( io_mem_0_r_bits_id ),
       .io_enq_bits_user( io_mem_0_r_bits_user ),
       .io_deq_ready( uncore_io_mem_0_r_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_resp( Queue_5_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_5_io_deq_bits_data ),
       .io_deq_bits_last( Queue_5_io_deq_bits_last ),
       .io_deq_bits_id( Queue_5_io_deq_bits_id ),
       .io_deq_bits_user( Queue_5_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( io_mem_0_b_valid ),
       .io_enq_bits_resp( io_mem_0_b_bits_resp ),
       .io_enq_bits_id( io_mem_0_b_bits_id ),
       .io_enq_bits_user( io_mem_0_b_bits_user ),
       .io_deq_ready( uncore_io_mem_0_b_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_resp( Queue_6_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_6_io_deq_bits_id ),
       .io_deq_bits_user( Queue_6_io_deq_bits_user )
       //.io_count(  )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T9(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

  reg [7:0] reg_R1A;
  reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
      reg_R1A = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge CLK) begin
    if (R1E) reg_R1A <= R1A;
    for (i = 0; i < 128; i=i+1) begin
      if (W0E && W0M[i]) ram[W0A][i] <= W0I[i];
    end
  end
  assign R1O = ram[reg_R1A];

endmodule

module MetadataArray_T6(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [87:0] W0I,
  input [87:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [87:0] R1O
);

  reg [5:0] reg_R1A;
  reg [87:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_R1A = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge CLK) begin
    if (R1E) reg_R1A <= R1A;
    for (i = 0; i < 88; i=i+1) begin
      if (W0E && W0M[i]) ram[W0A][i] <= W0I[i];
    end
  end
  assign R1O = ram[reg_R1A];

endmodule

module ICache_T178(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

  reg [7:0] reg_RW0A;
  reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
      reg_RW0A = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge CLK) begin
    if (RW0E && !RW0W) reg_RW0A <= RW0A;
    for (i = 0; i < 128; i=i+1) begin
      if (RW0E && RW0W) ram[RW0A][i] <= RW0I[i];
    end
  end
  assign RW0O = ram[reg_RW0A];

endmodule

module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [79:0] RW0M,
  input [79:0] RW0I,
  output [79:0] RW0O
);

  reg [5:0] reg_RW0A;
  reg [79:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0A = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge CLK) begin
    if (RW0E && !RW0W) reg_RW0A <= RW0A;
    for (i = 0; i < 80; i=i+1) begin
      if (RW0E && RW0W && RW0M[i]) ram[RW0A][i] <= RW0I[i];
    end
  end
  assign RW0O = ram[reg_RW0A];

endmodule


